magic
tech sky130A
timestamp 1697058477
<< nmos >>
rect 150 90 190 170
rect 250 90 290 170
<< ndiff >>
rect 95 150 150 170
rect 95 90 110 150
rect 130 90 150 150
rect 190 150 250 170
rect 190 90 210 150
rect 230 90 250 150
rect 290 150 370 170
rect 290 90 310 150
rect 330 90 370 150
rect 100 80 140 90
rect 200 80 240 90
rect 300 80 340 90
<< ndiffc >>
rect 110 90 130 150
rect 210 90 230 150
rect 310 90 330 150
<< psubdiff >>
rect 25 155 65 170
rect 25 110 35 155
rect 55 110 65 155
rect 25 90 65 110
<< psubdiffcont >>
rect 35 110 55 155
<< poly >>
rect 250 230 410 240
rect 0 220 190 230
rect 0 200 50 220
rect 70 200 190 220
rect 0 190 190 200
rect 150 170 190 190
rect 250 210 370 230
rect 390 210 410 230
rect 250 200 410 210
rect 250 170 290 200
rect 150 60 190 90
rect 250 60 290 90
<< polycont >>
rect 50 200 70 220
rect 370 210 390 230
<< locali >>
rect 300 380 340 410
rect 300 360 310 380
rect 330 360 340 380
rect 10 220 70 230
rect 10 200 20 220
rect 40 200 50 220
rect 10 190 70 200
rect 200 180 240 190
rect 20 155 70 170
rect 200 160 210 180
rect 230 160 240 180
rect 20 110 35 155
rect 55 110 70 155
rect 20 90 70 110
rect 20 65 30 90
rect 55 65 70 90
rect 20 60 70 65
rect 100 150 140 160
rect 100 90 110 150
rect 130 90 140 150
rect 100 70 140 90
rect 200 150 240 160
rect 200 90 210 150
rect 230 90 240 150
rect 200 80 240 90
rect 300 150 340 360
rect 360 230 410 240
rect 360 210 370 230
rect 390 210 410 230
rect 360 200 410 210
rect 300 90 310 150
rect 330 90 340 150
rect 300 80 340 90
rect 100 50 110 70
rect 130 50 140 70
rect 100 0 140 50
<< viali >>
rect 310 360 330 380
rect 20 200 40 220
rect 210 160 230 180
rect 30 65 55 90
rect 370 210 390 230
rect 110 50 130 70
<< metal1 >>
rect 300 640 350 650
rect 300 610 310 640
rect 340 610 350 640
rect 300 380 350 610
rect 300 360 310 380
rect 330 360 350 380
rect 300 350 350 360
rect 200 290 410 330
rect 0 220 50 230
rect 0 200 20 220
rect 40 200 50 220
rect 0 190 50 200
rect 200 180 240 290
rect 350 230 410 240
rect 350 210 370 230
rect 390 210 410 230
rect 350 200 410 210
rect 200 160 210 180
rect 230 160 240 180
rect 200 150 240 160
rect 20 90 70 110
rect 20 65 30 90
rect 55 65 70 90
rect 20 35 70 65
rect 20 5 30 35
rect 60 5 70 35
rect 20 0 70 5
rect 100 70 140 80
rect 100 50 110 70
rect 130 50 140 70
rect 100 35 140 50
rect 100 5 105 35
rect 135 5 140 35
rect 100 0 140 5
<< via1 >>
rect 310 610 340 640
rect 30 5 60 35
rect 105 5 135 35
<< metal2 >>
rect 0 640 350 650
rect 0 610 310 640
rect 340 610 350 640
rect 0 35 370 40
rect 0 5 30 35
rect 60 5 105 35
rect 135 5 370 35
rect 0 0 370 5
<< labels >>
rlabel metal2 0 610 10 650 3 VDD
port 1 e
rlabel metal2 0 0 10 40 3 VGND
port 2 e
rlabel metal1 0 190 20 230 1 VTAU
port 6 n
rlabel metal1 390 290 410 330 1 VOUT
port 7 n
rlabel metal1 400 200 410 240 7 VIN
port 8 w
<< end >>
