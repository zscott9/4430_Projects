magic
tech sky130A
timestamp 1695748008
<< nmos >>
rect 0 175 150 325
<< ndiff >>
rect -150 290 0 325
rect -150 210 -115 290
rect -35 210 0 290
rect -150 175 0 210
rect 150 290 300 325
rect 150 210 185 290
rect 265 210 300 290
rect 150 175 300 210
<< ndiffc >>
rect -115 210 -35 290
rect 185 210 265 290
<< psubdiff >>
rect -300 290 -150 325
rect -300 210 -265 290
rect -185 210 -150 290
rect -300 175 -150 210
<< psubdiffcont >>
rect -265 210 -185 290
<< poly >>
rect 0 325 150 500
rect 0 0 150 175
<< locali >>
rect -275 290 -25 300
rect -275 210 -265 290
rect -185 210 -115 290
rect -35 210 -25 290
rect -275 200 -25 210
rect 175 290 275 300
rect 175 210 185 290
rect 265 210 275 290
rect 175 200 275 210
<< end >>
