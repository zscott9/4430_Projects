magic
tech sky130A
timestamp 1697222590
<< nwell >>
rect 10 590 380 610
rect 10 460 600 590
rect 330 420 600 460
rect 330 410 590 420
rect 420 270 560 410
rect 420 240 790 270
rect 460 80 790 240
<< nmos >>
rect 280 290 320 370
rect 670 320 710 380
rect 180 100 220 180
rect 280 100 320 180
rect 870 70 930 450
<< pmos >>
rect 60 530 270 560
rect 380 480 430 570
rect 540 100 590 190
rect 640 100 690 190
<< ndiff >>
rect 840 420 870 450
rect 830 400 870 420
rect 230 360 280 370
rect 230 300 240 360
rect 270 300 280 360
rect 230 290 280 300
rect 320 360 360 370
rect 320 300 330 360
rect 350 300 360 360
rect 630 370 670 380
rect 630 330 640 370
rect 660 330 670 370
rect 630 320 670 330
rect 710 370 750 380
rect 710 330 720 370
rect 740 330 750 370
rect 710 320 750 330
rect 320 290 360 300
rect 140 170 180 180
rect 140 110 150 170
rect 170 110 180 170
rect 140 100 180 110
rect 220 170 280 180
rect 220 110 240 170
rect 270 110 280 170
rect 220 100 280 110
rect 320 160 360 180
rect 320 110 330 160
rect 350 130 360 160
rect 350 110 355 130
rect 320 100 355 110
rect 830 80 840 400
rect 860 80 870 400
rect 830 70 870 80
rect 930 420 960 450
rect 930 400 970 420
rect 930 80 940 400
rect 960 80 970 400
rect 930 70 970 80
<< pdiff >>
rect 60 585 270 590
rect 60 566 75 585
rect 250 566 270 585
rect 60 560 270 566
rect 340 560 380 570
rect 60 515 270 530
rect 60 490 70 515
rect 260 490 270 515
rect 60 485 270 490
rect 340 490 350 560
rect 370 490 380 560
rect 340 480 380 490
rect 430 550 510 570
rect 430 490 470 550
rect 500 490 510 550
rect 430 480 510 490
rect 490 170 540 190
rect 490 110 500 170
rect 530 110 540 170
rect 490 100 540 110
rect 590 180 640 190
rect 590 110 600 180
rect 630 110 640 180
rect 590 100 640 110
rect 690 180 760 190
rect 690 110 700 180
rect 730 110 760 180
rect 690 100 760 110
<< ndiffc >>
rect 240 300 270 360
rect 330 300 350 360
rect 640 330 660 370
rect 720 330 740 370
rect 150 110 170 170
rect 240 110 270 170
rect 330 110 350 160
rect 840 80 860 400
rect 940 80 960 400
<< pdiffc >>
rect 75 566 250 585
rect 70 490 260 515
rect 350 490 370 560
rect 470 490 500 550
rect 500 110 530 170
rect 600 110 630 180
rect 700 110 730 180
<< psubdiff >>
rect 50 240 100 260
rect 50 160 60 240
rect 90 160 100 240
rect 50 100 100 160
rect 385 80 440 100
rect 385 60 400 80
rect 420 60 440 80
rect 385 40 440 60
<< nsubdiff >>
rect 440 380 510 400
rect 440 340 460 380
rect 490 340 510 380
rect 440 320 510 340
<< psubdiffcont >>
rect 60 160 90 240
rect 400 60 420 80
<< nsubdiffcont >>
rect 460 340 490 380
<< poly >>
rect 290 580 430 600
rect 290 560 320 580
rect 380 570 430 580
rect 30 530 60 560
rect 270 530 320 560
rect 870 490 930 500
rect 380 450 430 480
rect 870 470 890 490
rect 920 470 930 490
rect 870 450 930 470
rect 200 430 320 440
rect 200 410 240 430
rect 270 410 320 430
rect 380 430 390 450
rect 420 430 430 450
rect 380 420 430 430
rect 670 440 720 450
rect 230 400 320 410
rect 670 410 680 440
rect 710 410 720 440
rect 670 400 720 410
rect 280 370 320 400
rect 670 380 710 400
rect 140 330 220 340
rect 140 300 150 330
rect 170 300 220 330
rect 140 290 220 300
rect 670 305 710 320
rect 180 180 220 290
rect 280 270 320 290
rect 540 270 690 280
rect 540 240 550 270
rect 580 240 690 270
rect 280 225 320 230
rect 280 220 325 225
rect 280 200 300 220
rect 320 200 325 220
rect 280 195 325 200
rect 540 220 690 240
rect 280 180 320 195
rect 540 190 590 220
rect 640 190 690 220
rect 180 40 220 100
rect 280 40 320 100
rect 540 60 590 100
rect 640 80 690 100
rect 870 40 930 70
<< polycont >>
rect 890 470 920 490
rect 240 410 270 430
rect 390 430 420 450
rect 680 410 710 440
rect 150 300 170 330
rect 550 240 580 270
rect 300 200 320 220
<< locali >>
rect 140 590 180 600
rect 60 585 150 590
rect 180 585 270 590
rect 60 566 75 585
rect 250 566 270 585
rect 760 570 800 580
rect 60 560 270 566
rect 340 560 380 570
rect 60 520 270 530
rect 60 515 160 520
rect 190 515 270 520
rect 60 490 70 515
rect 260 490 270 515
rect 60 485 270 490
rect 340 490 350 560
rect 370 490 380 560
rect 440 550 510 570
rect 760 560 770 570
rect 440 500 470 550
rect 340 480 380 490
rect 460 490 470 500
rect 500 490 510 550
rect 550 540 770 560
rect 800 540 990 560
rect 550 500 570 540
rect 460 480 510 490
rect 540 490 580 500
rect 330 450 430 480
rect 540 470 550 490
rect 570 470 580 490
rect 540 460 580 470
rect 720 490 930 500
rect 720 470 890 490
rect 920 470 930 490
rect 720 450 930 470
rect 200 430 280 440
rect 200 410 210 430
rect 230 410 240 430
rect 270 410 280 430
rect 330 430 390 450
rect 420 430 430 450
rect 330 420 430 430
rect 670 440 750 450
rect 220 360 280 380
rect 330 370 360 420
rect 670 410 680 440
rect 710 410 750 440
rect 970 420 990 540
rect 450 400 460 410
rect 70 330 180 340
rect 70 300 80 330
rect 110 300 150 330
rect 170 300 180 330
rect 70 290 180 300
rect 220 300 240 360
rect 270 300 280 360
rect 50 240 100 260
rect 50 160 60 240
rect 90 190 100 240
rect 90 170 180 190
rect 90 160 150 170
rect 50 140 150 160
rect 50 110 60 140
rect 90 110 150 140
rect 170 110 180 170
rect 50 90 180 110
rect 220 170 280 300
rect 320 360 360 370
rect 320 300 330 360
rect 350 300 360 360
rect 440 340 460 400
rect 490 340 510 410
rect 670 400 750 410
rect 440 320 510 340
rect 530 370 670 380
rect 530 360 640 370
rect 530 330 550 360
rect 570 330 640 360
rect 660 330 670 370
rect 530 320 670 330
rect 710 370 750 400
rect 710 330 720 370
rect 740 330 750 370
rect 320 290 360 300
rect 490 270 590 280
rect 490 240 550 270
rect 580 240 590 270
rect 300 220 360 230
rect 490 220 590 240
rect 710 270 750 330
rect 830 400 870 420
rect 320 200 360 220
rect 300 190 360 200
rect 490 170 540 220
rect 710 190 740 270
rect 220 110 240 170
rect 270 110 280 170
rect 220 90 280 110
rect 320 160 500 170
rect 320 110 330 160
rect 350 150 500 160
rect 350 130 360 150
rect 350 110 355 130
rect 320 100 355 110
rect 490 110 500 150
rect 530 110 540 170
rect 490 100 540 110
rect 590 180 640 190
rect 590 110 600 180
rect 630 110 640 180
rect 590 100 640 110
rect 690 180 740 190
rect 690 110 700 180
rect 730 110 740 180
rect 690 100 740 110
rect 390 80 430 90
rect 390 40 400 80
rect 420 60 430 80
rect 830 80 840 400
rect 860 80 870 400
rect 830 70 870 80
rect 930 400 990 420
rect 930 80 940 400
rect 960 350 990 400
rect 960 80 970 350
rect 930 70 970 80
<< viali >>
rect 150 585 180 590
rect 150 570 180 585
rect 160 515 190 520
rect 160 490 190 515
rect 470 520 500 540
rect 770 540 800 570
rect 550 470 570 490
rect 210 410 230 430
rect 80 300 110 330
rect 60 110 90 140
rect 460 380 490 410
rect 550 330 570 360
rect 360 200 380 220
rect 610 160 630 180
rect 840 80 860 100
rect 400 40 430 60
<< metal1 >>
rect 460 640 510 650
rect 140 610 150 640
rect 180 610 190 640
rect 140 590 190 610
rect 140 570 150 590
rect 180 570 190 590
rect 140 560 190 570
rect 460 610 470 640
rect 460 540 510 610
rect 150 520 200 530
rect 150 490 160 520
rect 190 490 200 520
rect 460 520 470 540
rect 500 520 510 540
rect 460 510 510 520
rect 620 640 660 650
rect 620 610 630 640
rect 150 480 200 490
rect 540 490 580 500
rect 540 480 550 490
rect 150 470 550 480
rect 570 470 580 490
rect 150 460 580 470
rect 620 460 660 610
rect 760 570 810 580
rect 760 540 770 570
rect 800 540 810 570
rect 760 510 810 540
rect 610 450 660 460
rect 180 430 240 440
rect 610 430 640 450
rect 180 410 210 430
rect 230 410 240 430
rect 180 400 240 410
rect 450 410 640 430
rect 450 380 460 410
rect 490 380 500 410
rect 450 370 500 380
rect 540 360 580 370
rect 30 330 120 340
rect 30 300 80 330
rect 110 300 120 330
rect 30 290 120 300
rect 540 330 550 360
rect 570 330 580 360
rect 340 220 440 230
rect 340 200 360 220
rect 380 200 440 220
rect 340 190 440 200
rect 50 140 100 160
rect 50 110 60 140
rect 90 110 100 140
rect 50 40 100 110
rect 50 10 60 40
rect 90 10 100 40
rect 50 0 100 10
rect 390 60 440 70
rect 390 40 400 60
rect 430 40 440 60
rect 390 30 440 40
rect 390 0 400 30
rect 430 0 440 30
rect 540 40 580 330
rect 610 190 640 410
rect 600 180 640 190
rect 600 160 610 180
rect 630 160 640 180
rect 600 150 640 160
rect 540 0 580 10
rect 830 100 870 110
rect 830 80 840 100
rect 860 80 870 100
rect 830 40 870 80
rect 830 0 870 10
<< via1 >>
rect 150 610 180 640
rect 470 610 510 640
rect 630 610 660 640
rect 60 10 90 40
rect 400 0 430 30
rect 540 10 580 40
rect 830 10 870 40
<< metal2 >>
rect 10 640 970 650
rect 10 610 150 640
rect 180 610 470 640
rect 510 610 630 640
rect 660 610 970 640
rect 0 10 60 40
rect 90 30 540 40
rect 90 10 400 30
rect 0 0 400 10
rect 430 10 540 30
rect 580 10 830 40
rect 870 10 970 40
rect 430 0 970 10
<< labels >>
rlabel metal1 30 290 50 340 1 VTAU
port 1 n
rlabel metal2 0 0 20 40 1 VGND
port 2 n
rlabel metal2 10 610 30 650 1 VDD
port 3 n
rlabel metal1 420 190 440 230 1 VIN2
port 5 n
rlabel metal1 180 400 200 440 1 VIN1
port 6 n
rlabel metal1 760 510 810 530 1 VOUT
port 7 n
rlabel locali 330 390 360 440 1 v34
rlabel locali 230 200 270 270 1 vint
rlabel locali 370 150 450 170 1 v56
rlabel locali 760 450 820 480 1 v78
<< end >>
