magic
tech sky130A
timestamp 1699640536
<< nmos >>
rect 0 0 90 90
<< ndiff >>
rect 0 -10 90 0
rect 0 -40 10 -10
rect 80 -40 90 -10
rect 0 -50 90 -40
<< ndiffc >>
rect 10 -40 80 -10
<< psubdiff >>
rect -160 80 -90 100
rect -160 50 -140 80
rect -110 50 -90 80
rect -160 30 -90 50
<< psubdiffcont >>
rect -140 50 -110 80
<< poly >>
rect -20 90 110 110
rect -20 0 0 90
rect 90 0 110 90
<< locali >>
rect -150 100 -100 120
rect -150 50 -140 100
rect -110 50 -100 100
rect -150 40 -100 50
rect 0 -10 90 0
rect 0 -40 10 -10
rect 80 -40 90 -10
rect 0 -50 90 -40
<< viali >>
rect -140 80 -110 100
rect 30 -40 60 -20
<< metal1 >>
rect -150 100 -100 140
rect -150 80 -140 100
rect -110 80 -100 100
rect -150 70 -100 80
rect 20 -20 70 -10
rect 20 -40 30 -20
rect 60 -40 70 -20
rect 20 -70 70 -40
<< labels >>
rlabel metal1 20 -70 70 -50 1 cap_in
port 1 n
rlabel metal1 -150 120 -100 140 1 GND
port 2 n
<< end >>
