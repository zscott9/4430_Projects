* NGSPICE file created from sky130_hilas_Bootstrap01.ext - technology: sky130A

.subckt sky130_hilas_Bootstrap01 RESIST VPWR VGND PBIAS NBIAS
X0 NBIAS PBIAS VPWR VPWR sky130_fd_pr__pfet_01v8 ad=1.68 pd=12.2 as=0.93 ps=6.13 w=5.81 l=0.2
X1 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X2 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X3 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X4 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X5 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=1.85 pd=12.5 as=0.924 ps=6.27 w=5.96 l=0.2
X6 VPWR PBIAS PBIAS VPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.13 as=1.74 ps=12.2 w=5.81 l=0.2
X7 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.983 ps=6.29 w=5.96 l=0.2
X8 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X9 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X10 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
R0 a_n535_n59# a_n454_n612# sky130_fd_pr__res_generic_po w=0.42 l=5.07
X11 NBIAS NBIAS VGND VGND sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.2
R1 a_n535_n59# RESIST sky130_fd_pr__res_generic_po w=0.42 l=5.07
X12 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X13 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X14 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X15 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.983 pd=6.29 as=1.73 ps=12.5 w=5.96 l=0.2
X16 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X17 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
X18 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0.924 pd=6.27 as=0.924 ps=6.27 w=5.96 l=0.2
.end

