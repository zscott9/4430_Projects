magic
tech sky130A
timestamp 1697207747
<< nmos >>
rect 280 290 320 370
rect 180 100 220 180
rect 280 100 320 180
<< ndiff >>
rect 230 360 280 370
rect 230 300 240 360
rect 270 300 280 360
rect 230 290 280 300
rect 320 360 360 370
rect 320 300 330 360
rect 350 300 360 360
rect 320 290 360 300
rect 140 170 180 180
rect 140 110 150 170
rect 170 110 180 170
rect 140 100 180 110
rect 220 170 280 180
rect 220 110 240 170
rect 270 110 280 170
rect 220 100 280 110
rect 320 160 360 180
rect 320 110 330 160
rect 350 110 360 160
rect 320 100 360 110
<< ndiffc >>
rect 240 300 270 360
rect 330 300 350 360
rect 150 110 170 170
rect 240 110 270 170
rect 330 110 350 160
<< psubdiff >>
rect 50 240 100 260
rect 50 160 60 240
rect 90 160 100 240
rect 50 100 100 160
<< psubdiffcont >>
rect 60 160 90 240
<< poly >>
rect 280 430 390 440
rect 280 400 350 430
rect 380 400 390 430
rect 280 390 390 400
rect 280 370 320 390
rect 140 330 220 340
rect 140 300 150 330
rect 170 300 220 330
rect 140 290 220 300
rect 180 180 220 290
rect 280 270 320 290
rect 280 220 360 230
rect 280 200 330 220
rect 350 200 360 220
rect 280 190 360 200
rect 280 180 320 190
rect 180 40 220 100
rect 280 40 320 100
<< polycont >>
rect 350 400 380 430
rect 150 300 170 330
rect 330 200 350 220
<< locali >>
rect 320 430 420 440
rect 320 400 350 430
rect 380 400 390 430
rect 410 400 420 430
rect 320 390 420 400
rect 220 360 280 380
rect 70 330 180 340
rect 70 300 80 330
rect 110 300 150 330
rect 170 300 180 330
rect 70 290 180 300
rect 220 300 240 360
rect 270 300 280 360
rect 50 240 100 260
rect 50 160 60 240
rect 90 190 100 240
rect 90 170 180 190
rect 90 160 150 170
rect 50 140 150 160
rect 50 110 60 140
rect 90 110 150 140
rect 170 110 180 170
rect 50 90 180 110
rect 220 170 280 300
rect 320 360 420 370
rect 320 300 330 360
rect 350 340 420 360
rect 350 320 390 340
rect 410 320 420 340
rect 350 300 420 320
rect 320 290 420 300
rect 320 220 360 230
rect 320 200 330 220
rect 350 200 360 220
rect 320 190 360 200
rect 220 110 240 170
rect 270 110 280 170
rect 220 90 280 110
rect 320 160 390 170
rect 320 110 330 160
rect 350 150 390 160
rect 350 120 370 150
rect 350 110 390 120
rect 320 100 390 110
<< viali >>
rect 390 400 410 430
rect 80 300 110 330
rect 60 110 90 140
rect 390 320 410 340
rect 360 200 380 220
rect 370 120 390 150
<< metal1 >>
rect 460 640 500 650
rect 460 610 470 640
rect 340 430 440 440
rect 340 400 390 430
rect 410 400 440 430
rect 340 390 440 400
rect 460 350 500 610
rect 380 340 500 350
rect 30 330 120 340
rect 30 300 80 330
rect 110 300 120 330
rect 380 320 390 340
rect 410 320 500 340
rect 380 310 500 320
rect 30 290 120 300
rect 320 220 440 230
rect 320 200 360 220
rect 380 200 440 220
rect 320 190 440 200
rect 460 160 500 310
rect 50 140 100 160
rect 50 110 60 140
rect 90 110 100 140
rect 360 150 500 160
rect 360 120 370 150
rect 390 120 500 150
rect 360 110 500 120
rect 50 40 100 110
rect 50 10 60 40
rect 90 10 100 40
rect 50 0 100 10
<< via1 >>
rect 470 610 500 640
rect 60 10 90 40
<< metal2 >>
rect 10 640 510 650
rect 10 610 470 640
rect 500 610 510 640
rect 0 10 60 40
rect 90 10 510 40
rect 0 0 510 10
<< labels >>
rlabel metal1 30 290 50 340 1 VTAU
port 1 n
rlabel metal2 0 0 20 40 1 VGND
port 2 n
rlabel metal2 10 610 30 650 1 VDD
port 3 n
rlabel metal1 420 390 440 440 1 VIN1
port 4 n
rlabel metal1 420 190 440 230 1 VIN2
port 5 n
<< end >>
