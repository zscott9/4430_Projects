magic
tech sky130A
timestamp 1697480338
<< nwell >>
rect 0 210 520 590
rect 0 50 1020 210
<< nmos >>
rect 610 450 650 530
rect 790 439 830 530
rect 610 280 650 360
rect 790 280 830 360
rect 880 280 920 360
<< pmos >>
rect 90 80 130 240
rect 270 80 310 560
rect 360 80 400 560
<< ndiff >>
rect 560 520 610 530
rect 560 460 570 520
rect 600 460 610 520
rect 560 450 610 460
rect 650 450 700 530
rect 740 520 790 530
rect 740 450 750 520
rect 780 450 790 520
rect 740 439 790 450
rect 830 439 880 530
rect 560 350 610 360
rect 560 290 570 350
rect 600 290 610 350
rect 560 280 610 290
rect 650 280 700 360
rect 740 350 790 360
rect 740 290 750 350
rect 780 290 790 350
rect 740 280 790 290
rect 830 350 880 360
rect 830 290 840 350
rect 870 290 880 350
rect 830 280 880 290
rect 920 280 970 360
<< pdiff >>
rect 220 550 270 560
rect 40 230 90 240
rect 40 90 50 230
rect 80 90 90 230
rect 40 80 90 90
rect 130 230 180 240
rect 130 90 140 230
rect 170 90 180 230
rect 130 80 180 90
rect 220 90 230 550
rect 260 90 270 550
rect 220 80 270 90
rect 310 550 360 560
rect 310 90 320 550
rect 350 90 360 550
rect 310 80 360 90
rect 400 550 450 560
rect 400 90 410 550
rect 440 90 450 550
rect 400 80 450 90
<< ndiffc >>
rect 570 460 600 520
rect 750 450 780 520
rect 570 290 600 350
rect 750 290 780 350
rect 840 290 870 350
<< pdiffc >>
rect 50 90 80 230
rect 140 90 170 230
rect 230 90 260 550
rect 320 90 350 550
rect 410 90 440 550
<< nsubdiff >>
rect 40 530 170 570
rect 40 400 80 530
rect 130 400 170 530
rect 40 360 170 400
<< nsubdiffcont >>
rect 80 400 130 530
<< poly >>
rect 270 610 310 620
rect 270 590 280 610
rect 300 590 310 610
rect 270 560 310 590
rect 360 610 400 620
rect 360 590 370 610
rect 390 590 400 610
rect 360 560 400 590
rect 610 580 650 590
rect 610 560 620 580
rect 640 560 650 580
rect 90 290 130 300
rect 90 270 100 290
rect 120 270 130 290
rect 90 240 130 270
rect 610 530 650 560
rect 790 530 830 550
rect 610 360 650 450
rect 790 420 830 439
rect 790 360 830 380
rect 880 360 920 380
rect 610 250 650 280
rect 790 250 830 280
rect 790 230 800 250
rect 820 230 830 250
rect 790 220 830 230
rect 880 250 920 280
rect 880 230 890 250
rect 910 230 920 250
rect 880 220 920 230
rect 90 60 130 80
rect 270 60 310 80
rect 360 60 400 80
<< polycont >>
rect 280 590 300 610
rect 370 590 390 610
rect 620 560 640 580
rect 100 270 120 290
rect 800 230 820 250
rect 890 230 910 250
<< locali >>
rect 270 610 310 620
rect 270 590 280 610
rect 300 590 310 610
rect 270 580 310 590
rect 360 610 400 620
rect 360 590 370 610
rect 390 590 400 610
rect 360 580 400 590
rect 610 580 650 590
rect 570 560 620 580
rect 640 560 650 580
rect 220 550 270 560
rect 70 530 90 550
rect 120 530 140 550
rect 70 400 80 530
rect 130 400 140 530
rect 70 390 140 400
rect 90 290 130 300
rect 90 270 100 290
rect 120 270 130 290
rect 90 260 130 270
rect 40 230 90 240
rect 40 90 50 230
rect 80 90 90 230
rect 40 80 90 90
rect 130 230 180 240
rect 130 90 140 230
rect 170 90 180 230
rect 130 80 180 90
rect 220 90 230 550
rect 260 90 270 550
rect 220 80 270 90
rect 310 550 360 560
rect 310 90 320 550
rect 350 90 360 550
rect 310 80 360 90
rect 400 550 450 560
rect 400 90 410 550
rect 440 90 450 550
rect 570 550 650 560
rect 570 530 600 550
rect 560 520 610 530
rect 560 460 570 520
rect 600 460 610 520
rect 560 450 610 460
rect 650 450 700 530
rect 740 520 790 530
rect 740 450 750 520
rect 780 450 790 520
rect 660 360 690 450
rect 740 439 790 450
rect 560 350 610 360
rect 560 290 570 350
rect 600 290 610 350
rect 560 280 610 290
rect 650 320 700 360
rect 650 290 660 320
rect 690 290 700 320
rect 650 280 700 290
rect 740 350 790 360
rect 740 290 750 350
rect 780 290 790 350
rect 740 260 790 290
rect 830 350 880 360
rect 830 290 840 350
rect 870 290 880 350
rect 830 280 880 290
rect 740 230 750 260
rect 780 250 920 260
rect 780 230 800 250
rect 820 230 890 250
rect 910 230 920 250
rect 740 220 920 230
rect 400 80 450 90
<< viali >>
rect 280 590 300 610
rect 370 590 390 610
rect 90 530 120 550
rect 100 270 120 290
rect 50 140 80 170
rect 140 90 170 120
rect 230 480 260 510
rect 320 90 350 120
rect 410 180 440 210
rect 570 480 600 510
rect 750 450 780 480
rect 570 320 600 350
rect 660 290 690 320
rect 840 290 870 320
rect 750 230 780 260
<< metal1 >>
rect 80 610 90 640
rect 120 610 130 640
rect 270 610 310 620
rect 360 610 400 620
rect 80 550 130 610
rect 240 590 280 610
rect 300 590 310 610
rect 330 590 370 610
rect 390 590 400 610
rect 270 580 310 590
rect 360 580 400 590
rect 80 530 90 550
rect 120 530 130 550
rect 80 520 130 530
rect 220 510 610 520
rect 220 480 230 510
rect 260 480 570 510
rect 600 480 610 510
rect 220 470 610 480
rect 740 480 790 490
rect 740 450 750 480
rect 780 450 790 480
rect 740 420 790 450
rect 560 380 790 420
rect 560 350 610 380
rect 560 320 570 350
rect 600 320 610 350
rect 560 310 610 320
rect 650 320 700 330
rect 50 290 130 300
rect 50 270 100 290
rect 120 270 130 290
rect 50 260 130 270
rect 650 290 660 320
rect 690 290 700 320
rect 400 210 450 220
rect 400 180 410 210
rect 440 180 450 210
rect 40 170 90 180
rect 400 170 450 180
rect 40 140 50 170
rect 80 140 90 170
rect 40 130 90 140
rect 130 120 360 130
rect 130 90 140 120
rect 170 90 320 120
rect 350 90 360 120
rect 130 80 360 90
rect 650 40 700 290
rect 830 320 880 330
rect 830 290 840 320
rect 870 290 880 320
rect 740 260 790 270
rect 740 230 750 260
rect 780 230 790 260
rect 740 210 790 230
rect 740 180 750 210
rect 780 180 790 210
rect 740 170 790 180
rect 650 10 660 40
rect 690 10 700 40
rect 650 0 700 10
rect 830 40 880 290
rect 830 10 840 40
rect 870 10 880 40
rect 830 0 880 10
<< via1 >>
rect 90 610 120 640
rect 410 180 440 210
rect 50 140 80 170
rect 750 180 780 210
rect 660 10 690 40
rect 840 10 870 40
<< metal2 >>
rect 0 640 1760 650
rect 0 610 90 640
rect 120 610 1760 640
rect 50 180 80 610
rect 400 210 790 220
rect 400 180 410 210
rect 440 180 750 210
rect 780 180 790 210
rect 40 170 90 180
rect 400 170 790 180
rect 40 140 50 170
rect 80 140 90 170
rect 40 130 90 140
rect 0 10 660 40
rect 690 10 840 40
rect 870 10 1760 40
rect 0 0 1760 10
<< labels >>
rlabel metal1 50 260 70 300 1 VTAU
port 1 n
rlabel metal2 0 610 20 650 1 VDD
port 2 n
rlabel metal1 240 590 260 610 1 VIN1
port 3 n
rlabel metal1 330 590 350 610 1 VIN2
port 4 n
rlabel metal1 520 470 560 520 1 v13
rlabel metal2 0 0 20 40 1 VGND
port 5 n
rlabel metal2 520 170 600 220 1 V26
rlabel metal1 740 380 790 420 1 V45
<< end >>
