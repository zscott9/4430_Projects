magic
tech sky130A
timestamp 1702459089
<< nwell >>
rect 2720 1940 3020 1980
rect 5740 1940 6080 1980
rect 2010 1750 2580 1940
rect 2720 1750 4190 1940
rect 5030 1750 5600 1940
rect 5740 1750 7200 1940
rect 2720 1460 3020 1750
rect 5740 1460 6040 1750
rect 7470 1410 7790 1980
rect 8800 1910 9140 1990
rect 8490 1580 9140 1910
rect 10010 1770 10580 1960
rect 11050 1770 12190 1960
rect 7920 1410 8180 1550
rect 8800 1420 9140 1580
rect 7920 1400 8090 1410
<< nmos >>
rect 1210 1500 1910 1980
rect 2100 1530 2140 1670
rect 2380 1530 2420 1670
rect 3130 1530 3170 1670
rect 3420 1530 3460 1670
rect 3700 1530 3740 1670
rect 3990 1530 4030 1670
rect 4270 1500 4970 1980
rect 5120 1530 5160 1670
rect 5400 1530 5440 1670
rect 2590 1450 2680 1470
rect 7330 1750 7370 1830
rect 6150 1530 6190 1670
rect 6430 1530 6470 1670
rect 6720 1530 6760 1670
rect 7000 1530 7040 1670
rect 7330 1610 7370 1690
rect 5610 1450 5700 1470
rect 8010 1640 8050 1820
rect 8330 1610 8370 1850
rect 9210 1520 9910 2000
rect 10100 1550 10140 1690
rect 10380 1550 10420 1690
rect 10880 1500 10920 1980
rect 11140 1550 11180 1690
rect 11420 1550 11460 1690
rect 11700 1550 11740 1690
rect 11990 1550 12030 1690
rect 10610 1470 10700 1490
<< pmos >>
rect 2100 1780 2140 1920
rect 2380 1780 2420 1920
rect 2880 1480 2920 1960
rect 3130 1780 3170 1920
rect 3420 1780 3460 1920
rect 3700 1780 3740 1920
rect 3990 1780 4030 1920
rect 5120 1780 5160 1920
rect 5400 1780 5440 1920
rect 5900 1480 5940 1960
rect 6150 1780 6190 1920
rect 6430 1780 6470 1920
rect 6720 1780 6760 1920
rect 7000 1780 7040 1920
rect 7640 1440 7680 1920
rect 8690 1610 8730 1850
rect 8060 1460 8100 1500
rect 8980 1450 9020 1930
rect 10100 1800 10140 1940
rect 10380 1800 10420 1940
rect 11140 1800 11180 1940
rect 11420 1800 11460 1940
rect 11700 1800 11740 1940
rect 11990 1800 12030 1940
<< ndiff >>
rect 2030 1650 2100 1670
rect 2030 1550 2050 1650
rect 2080 1550 2100 1650
rect 2030 1530 2100 1550
rect 2140 1650 2210 1670
rect 2140 1550 2160 1650
rect 2190 1550 2210 1650
rect 2140 1530 2210 1550
rect 2310 1650 2380 1670
rect 2310 1550 2330 1650
rect 2360 1550 2380 1650
rect 2310 1530 2380 1550
rect 2420 1650 2490 1670
rect 2420 1550 2440 1650
rect 2470 1550 2490 1650
rect 2420 1530 2490 1550
rect 2590 1600 2680 1610
rect 2590 1580 2620 1600
rect 2640 1580 2680 1600
rect 1210 1470 1910 1500
rect 2590 1470 2680 1580
rect 3060 1650 3130 1670
rect 3060 1550 3080 1650
rect 3110 1550 3130 1650
rect 3060 1530 3130 1550
rect 3170 1650 3240 1670
rect 3170 1550 3190 1650
rect 3220 1550 3240 1650
rect 3170 1530 3240 1550
rect 3350 1650 3420 1670
rect 3350 1550 3370 1650
rect 3400 1550 3420 1650
rect 3350 1530 3420 1550
rect 3460 1650 3530 1670
rect 3460 1550 3480 1650
rect 3510 1550 3530 1650
rect 3460 1530 3530 1550
rect 3630 1650 3700 1670
rect 3630 1550 3650 1650
rect 3680 1550 3700 1650
rect 3630 1530 3700 1550
rect 3740 1650 3810 1670
rect 3740 1550 3760 1650
rect 3790 1550 3810 1650
rect 3740 1530 3810 1550
rect 3920 1650 3990 1670
rect 3920 1550 3940 1650
rect 3970 1550 3990 1650
rect 3920 1530 3990 1550
rect 4030 1650 4100 1670
rect 4030 1550 4050 1650
rect 4080 1550 4100 1650
rect 4030 1530 4100 1550
rect 5050 1650 5120 1670
rect 5050 1550 5070 1650
rect 5100 1550 5120 1650
rect 5050 1530 5120 1550
rect 5160 1650 5230 1670
rect 5160 1550 5180 1650
rect 5210 1550 5230 1650
rect 5160 1530 5230 1550
rect 5330 1650 5400 1670
rect 5330 1550 5350 1650
rect 5380 1550 5400 1650
rect 5330 1530 5400 1550
rect 5440 1650 5510 1670
rect 5440 1550 5460 1650
rect 5490 1550 5510 1650
rect 5440 1530 5510 1550
rect 5610 1600 5700 1610
rect 5610 1580 5650 1600
rect 5670 1580 5700 1600
rect 1210 1430 1670 1470
rect 1730 1430 1810 1470
rect 1870 1430 1910 1470
rect 1210 1400 1910 1430
rect 2590 1420 2680 1450
rect 4270 1470 4970 1500
rect 5610 1470 5700 1580
rect 7280 1810 7330 1830
rect 7280 1770 7300 1810
rect 7320 1770 7330 1810
rect 7280 1750 7330 1770
rect 7370 1810 7430 1830
rect 7370 1770 7390 1810
rect 7410 1770 7430 1810
rect 7370 1750 7430 1770
rect 7280 1670 7330 1690
rect 6080 1650 6150 1670
rect 6080 1550 6100 1650
rect 6130 1550 6150 1650
rect 6080 1530 6150 1550
rect 6190 1650 6260 1670
rect 6190 1550 6210 1650
rect 6240 1550 6260 1650
rect 6190 1530 6260 1550
rect 6360 1650 6430 1670
rect 6360 1550 6380 1650
rect 6410 1550 6430 1650
rect 6360 1530 6430 1550
rect 6470 1650 6540 1670
rect 6470 1550 6490 1650
rect 6520 1550 6540 1650
rect 6470 1530 6540 1550
rect 6650 1650 6720 1670
rect 6650 1550 6670 1650
rect 6700 1550 6720 1650
rect 6650 1530 6720 1550
rect 6760 1650 6830 1670
rect 6760 1550 6780 1650
rect 6810 1550 6830 1650
rect 6760 1530 6830 1550
rect 6930 1650 7000 1670
rect 6930 1550 6950 1650
rect 6980 1550 7000 1650
rect 6930 1530 7000 1550
rect 7040 1650 7110 1670
rect 7040 1550 7060 1650
rect 7090 1550 7110 1650
rect 7280 1630 7300 1670
rect 7320 1630 7330 1670
rect 7280 1610 7330 1630
rect 7370 1670 7430 1690
rect 7370 1630 7390 1670
rect 7410 1630 7430 1670
rect 7370 1610 7430 1630
rect 7040 1530 7110 1550
rect 4270 1440 4730 1470
rect 4790 1440 4870 1470
rect 4930 1440 4970 1470
rect 4270 1430 4970 1440
rect 5610 1420 5700 1450
rect 8250 1830 8330 1850
rect 7920 1800 8010 1820
rect 7920 1660 7940 1800
rect 7990 1660 8010 1800
rect 7920 1640 8010 1660
rect 8050 1800 8140 1820
rect 8050 1660 8070 1800
rect 8120 1660 8140 1800
rect 8050 1640 8140 1660
rect 8250 1630 8270 1830
rect 8310 1630 8330 1830
rect 8250 1610 8330 1630
rect 8370 1830 8450 1850
rect 8370 1630 8390 1830
rect 8430 1630 8450 1830
rect 8370 1610 8450 1630
rect 10800 1950 10880 1980
rect 10030 1670 10100 1690
rect 10030 1570 10050 1670
rect 10080 1570 10100 1670
rect 10030 1550 10100 1570
rect 10140 1670 10210 1690
rect 10140 1570 10160 1670
rect 10190 1570 10210 1670
rect 10140 1550 10210 1570
rect 10310 1670 10380 1690
rect 10310 1570 10330 1670
rect 10360 1570 10380 1670
rect 10310 1550 10380 1570
rect 10420 1670 10490 1690
rect 10420 1570 10440 1670
rect 10470 1570 10490 1670
rect 10420 1550 10490 1570
rect 10610 1610 10700 1630
rect 10610 1590 10650 1610
rect 10670 1590 10700 1610
rect 9210 1490 9910 1520
rect 10610 1490 10700 1590
rect 10800 1530 10830 1950
rect 10850 1530 10880 1950
rect 10800 1500 10880 1530
rect 10920 1950 11000 1980
rect 10920 1530 10950 1950
rect 10970 1530 11000 1950
rect 11070 1670 11140 1690
rect 11070 1570 11090 1670
rect 11120 1570 11140 1670
rect 11070 1550 11140 1570
rect 11180 1670 11250 1690
rect 11180 1570 11200 1670
rect 11230 1570 11250 1670
rect 11180 1550 11250 1570
rect 11350 1670 11420 1690
rect 11350 1570 11370 1670
rect 11400 1570 11420 1670
rect 11350 1550 11420 1570
rect 11460 1670 11530 1690
rect 11460 1570 11480 1670
rect 11510 1570 11530 1670
rect 11460 1550 11530 1570
rect 11630 1670 11700 1690
rect 11630 1570 11650 1670
rect 11680 1570 11700 1670
rect 11630 1550 11700 1570
rect 11740 1670 11810 1690
rect 11740 1570 11760 1670
rect 11790 1570 11810 1670
rect 11740 1550 11810 1570
rect 11920 1670 11990 1690
rect 11920 1570 11940 1670
rect 11970 1570 11990 1670
rect 11920 1550 11990 1570
rect 12030 1670 12100 1690
rect 12030 1570 12050 1670
rect 12080 1570 12100 1670
rect 12030 1550 12100 1570
rect 10920 1500 11000 1530
rect 9210 1450 9670 1490
rect 9730 1450 9810 1490
rect 9870 1450 9910 1490
rect 9210 1420 9910 1450
rect 10610 1440 10700 1470
<< pdiff >>
rect 2800 1930 2880 1960
rect 2030 1900 2100 1920
rect 2030 1800 2050 1900
rect 2080 1800 2100 1900
rect 2030 1780 2100 1800
rect 2140 1900 2210 1920
rect 2140 1800 2160 1900
rect 2190 1800 2210 1900
rect 2140 1780 2210 1800
rect 2310 1900 2380 1920
rect 2310 1800 2330 1900
rect 2360 1800 2380 1900
rect 2310 1780 2380 1800
rect 2420 1900 2490 1920
rect 2420 1800 2440 1900
rect 2470 1800 2490 1900
rect 2420 1780 2490 1800
rect 2800 1510 2830 1930
rect 2850 1510 2880 1930
rect 2800 1480 2880 1510
rect 2920 1930 3000 1960
rect 2920 1510 2950 1930
rect 2970 1510 3000 1930
rect 3060 1900 3130 1920
rect 3060 1800 3080 1900
rect 3110 1800 3130 1900
rect 3060 1780 3130 1800
rect 3170 1900 3240 1920
rect 3170 1800 3190 1900
rect 3220 1800 3240 1900
rect 3170 1780 3240 1800
rect 3350 1900 3420 1920
rect 3350 1800 3370 1900
rect 3400 1800 3420 1900
rect 3350 1780 3420 1800
rect 3460 1900 3530 1920
rect 3460 1800 3480 1900
rect 3510 1800 3530 1900
rect 3460 1780 3530 1800
rect 3630 1900 3700 1920
rect 3630 1800 3650 1900
rect 3680 1800 3700 1900
rect 3630 1780 3700 1800
rect 3740 1900 3810 1920
rect 3740 1800 3760 1900
rect 3790 1800 3810 1900
rect 3740 1780 3810 1800
rect 3920 1900 3990 1920
rect 3920 1800 3940 1900
rect 3970 1800 3990 1900
rect 3920 1780 3990 1800
rect 4030 1900 4100 1920
rect 4030 1800 4050 1900
rect 4080 1800 4100 1900
rect 4030 1780 4100 1800
rect 2920 1480 3000 1510
rect 5820 1930 5900 1960
rect 5050 1900 5120 1920
rect 5050 1800 5070 1900
rect 5100 1800 5120 1900
rect 5050 1780 5120 1800
rect 5160 1900 5230 1920
rect 5160 1800 5180 1900
rect 5210 1800 5230 1900
rect 5160 1780 5230 1800
rect 5330 1900 5400 1920
rect 5330 1800 5350 1900
rect 5380 1800 5400 1900
rect 5330 1780 5400 1800
rect 5440 1900 5510 1920
rect 5440 1800 5460 1900
rect 5490 1800 5510 1900
rect 5440 1780 5510 1800
rect 5820 1510 5850 1930
rect 5870 1510 5900 1930
rect 5820 1480 5900 1510
rect 5940 1930 6020 1960
rect 5940 1510 5970 1930
rect 5990 1510 6020 1930
rect 6080 1900 6150 1920
rect 6080 1800 6100 1900
rect 6130 1800 6150 1900
rect 6080 1780 6150 1800
rect 6190 1900 6260 1920
rect 6190 1800 6210 1900
rect 6240 1800 6260 1900
rect 6190 1780 6260 1800
rect 6360 1900 6430 1920
rect 6360 1800 6380 1900
rect 6410 1800 6430 1900
rect 6360 1780 6430 1800
rect 6470 1900 6540 1920
rect 6470 1800 6490 1900
rect 6520 1800 6540 1900
rect 6470 1780 6540 1800
rect 6650 1900 6720 1920
rect 6650 1800 6670 1900
rect 6700 1800 6720 1900
rect 6650 1780 6720 1800
rect 6760 1900 6830 1920
rect 6760 1800 6780 1900
rect 6810 1800 6830 1900
rect 6760 1780 6830 1800
rect 6930 1900 7000 1920
rect 6930 1800 6950 1900
rect 6980 1800 7000 1900
rect 6930 1780 7000 1800
rect 7040 1900 7110 1920
rect 7040 1800 7060 1900
rect 7090 1800 7110 1900
rect 7560 1890 7640 1920
rect 7040 1780 7110 1800
rect 5940 1480 6020 1510
rect 7560 1470 7590 1890
rect 7610 1470 7640 1890
rect 7560 1440 7640 1470
rect 7680 1890 7760 1920
rect 7680 1470 7710 1890
rect 7730 1470 7760 1890
rect 8900 1900 8980 1930
rect 8610 1830 8690 1850
rect 8610 1630 8630 1830
rect 8670 1630 8690 1830
rect 8610 1610 8690 1630
rect 8730 1830 8810 1850
rect 8730 1630 8750 1830
rect 8790 1630 8810 1830
rect 8730 1610 8810 1630
rect 7680 1440 7760 1470
rect 8000 1490 8060 1500
rect 8000 1470 8020 1490
rect 8040 1470 8060 1490
rect 8000 1460 8060 1470
rect 8100 1490 8160 1500
rect 8100 1470 8120 1490
rect 8140 1470 8160 1490
rect 8100 1460 8160 1470
rect 8900 1480 8930 1900
rect 8950 1480 8980 1900
rect 8900 1450 8980 1480
rect 9020 1900 9100 1930
rect 9020 1480 9050 1900
rect 9070 1480 9100 1900
rect 10030 1920 10100 1940
rect 10030 1820 10050 1920
rect 10080 1820 10100 1920
rect 10030 1800 10100 1820
rect 10140 1920 10210 1940
rect 10140 1820 10160 1920
rect 10190 1820 10210 1920
rect 10140 1800 10210 1820
rect 10310 1920 10380 1940
rect 10310 1820 10330 1920
rect 10360 1820 10380 1920
rect 10310 1800 10380 1820
rect 10420 1920 10490 1940
rect 10420 1820 10440 1920
rect 10470 1820 10490 1920
rect 10420 1800 10490 1820
rect 9020 1450 9100 1480
rect 11070 1920 11140 1940
rect 11070 1820 11090 1920
rect 11120 1820 11140 1920
rect 11070 1800 11140 1820
rect 11180 1920 11250 1940
rect 11180 1820 11200 1920
rect 11230 1820 11250 1920
rect 11180 1800 11250 1820
rect 11350 1920 11420 1940
rect 11350 1820 11370 1920
rect 11400 1820 11420 1920
rect 11350 1800 11420 1820
rect 11460 1920 11530 1940
rect 11460 1820 11480 1920
rect 11510 1820 11530 1920
rect 11460 1800 11530 1820
rect 11630 1920 11700 1940
rect 11630 1820 11650 1920
rect 11680 1820 11700 1920
rect 11630 1800 11700 1820
rect 11740 1920 11810 1940
rect 11740 1820 11760 1920
rect 11790 1820 11810 1920
rect 11740 1800 11810 1820
rect 11920 1920 11990 1940
rect 11920 1820 11940 1920
rect 11970 1820 11990 1920
rect 11920 1800 11990 1820
rect 12030 1920 12100 1940
rect 12030 1820 12050 1920
rect 12080 1820 12100 1920
rect 12030 1800 12100 1820
<< ndiffc >>
rect 2050 1550 2080 1650
rect 2160 1550 2190 1650
rect 2330 1550 2360 1650
rect 2440 1550 2470 1650
rect 2620 1580 2640 1600
rect 3080 1550 3110 1650
rect 3190 1550 3220 1650
rect 3370 1550 3400 1650
rect 3480 1550 3510 1650
rect 3650 1550 3680 1650
rect 3760 1550 3790 1650
rect 3940 1550 3970 1650
rect 4050 1550 4080 1650
rect 5070 1550 5100 1650
rect 5180 1550 5210 1650
rect 5350 1550 5380 1650
rect 5460 1550 5490 1650
rect 5650 1580 5670 1600
rect 1670 1430 1730 1470
rect 1810 1430 1870 1470
rect 7300 1770 7320 1810
rect 7390 1770 7410 1810
rect 6100 1550 6130 1650
rect 6210 1550 6240 1650
rect 6380 1550 6410 1650
rect 6490 1550 6520 1650
rect 6670 1550 6700 1650
rect 6780 1550 6810 1650
rect 6950 1550 6980 1650
rect 7060 1550 7090 1650
rect 7300 1630 7320 1670
rect 7390 1630 7410 1670
rect 4730 1440 4790 1470
rect 4870 1440 4930 1470
rect 7940 1660 7990 1800
rect 8070 1660 8120 1800
rect 8270 1630 8310 1830
rect 8390 1630 8430 1830
rect 10050 1570 10080 1670
rect 10160 1570 10190 1670
rect 10330 1570 10360 1670
rect 10440 1570 10470 1670
rect 10650 1590 10670 1610
rect 10830 1530 10850 1950
rect 10950 1530 10970 1950
rect 11090 1570 11120 1670
rect 11200 1570 11230 1670
rect 11370 1570 11400 1670
rect 11480 1570 11510 1670
rect 11650 1570 11680 1670
rect 11760 1570 11790 1670
rect 11940 1570 11970 1670
rect 12050 1570 12080 1670
rect 9670 1450 9730 1490
rect 9810 1450 9870 1490
<< pdiffc >>
rect 2050 1800 2080 1900
rect 2160 1800 2190 1900
rect 2330 1800 2360 1900
rect 2440 1800 2470 1900
rect 2830 1510 2850 1930
rect 2950 1510 2970 1930
rect 3080 1800 3110 1900
rect 3190 1800 3220 1900
rect 3370 1800 3400 1900
rect 3480 1800 3510 1900
rect 3650 1800 3680 1900
rect 3760 1800 3790 1900
rect 3940 1800 3970 1900
rect 4050 1800 4080 1900
rect 5070 1800 5100 1900
rect 5180 1800 5210 1900
rect 5350 1800 5380 1900
rect 5460 1800 5490 1900
rect 5850 1510 5870 1930
rect 5970 1510 5990 1930
rect 6100 1800 6130 1900
rect 6210 1800 6240 1900
rect 6380 1800 6410 1900
rect 6490 1800 6520 1900
rect 6670 1800 6700 1900
rect 6780 1800 6810 1900
rect 6950 1800 6980 1900
rect 7060 1800 7090 1900
rect 7590 1470 7610 1890
rect 7710 1470 7730 1890
rect 8630 1630 8670 1830
rect 8750 1630 8790 1830
rect 8020 1470 8040 1490
rect 8120 1470 8140 1490
rect 8930 1480 8950 1900
rect 9050 1480 9070 1900
rect 10050 1820 10080 1920
rect 10160 1820 10190 1920
rect 10330 1820 10360 1920
rect 10440 1820 10470 1920
rect 11090 1820 11120 1920
rect 11200 1820 11230 1920
rect 11370 1820 11400 1920
rect 11480 1820 11510 1920
rect 11650 1820 11680 1920
rect 11760 1820 11790 1920
rect 11940 1820 11970 1920
rect 12050 1820 12080 1920
<< psubdiff >>
rect 2210 1650 2280 1670
rect 2210 1550 2230 1650
rect 2260 1550 2280 1650
rect 2210 1530 2280 1550
rect 2490 1650 2560 1670
rect 2490 1550 2510 1650
rect 2540 1550 2560 1650
rect 2490 1530 2560 1550
rect 3240 1650 3310 1670
rect 3240 1550 3260 1650
rect 3290 1550 3310 1650
rect 3240 1530 3310 1550
rect 3530 1650 3600 1670
rect 3530 1550 3550 1650
rect 3580 1550 3600 1650
rect 3530 1530 3600 1550
rect 3810 1650 3880 1670
rect 3810 1550 3830 1650
rect 3860 1550 3880 1650
rect 3810 1530 3880 1550
rect 4100 1650 4170 1670
rect 4100 1550 4120 1650
rect 4150 1550 4170 1650
rect 4100 1530 4170 1550
rect 5230 1650 5300 1670
rect 5230 1550 5250 1650
rect 5280 1550 5300 1650
rect 5230 1530 5300 1550
rect 5510 1650 5580 1670
rect 5510 1550 5530 1650
rect 5560 1550 5580 1650
rect 5510 1530 5580 1550
rect 7220 1810 7280 1830
rect 7220 1770 7240 1810
rect 7260 1770 7280 1810
rect 7220 1750 7280 1770
rect 7220 1670 7280 1690
rect 6260 1650 6330 1670
rect 6260 1550 6280 1650
rect 6310 1550 6330 1650
rect 6260 1530 6330 1550
rect 6540 1650 6610 1670
rect 6540 1550 6560 1650
rect 6590 1550 6610 1650
rect 6540 1530 6610 1550
rect 6830 1650 6900 1670
rect 6830 1550 6850 1650
rect 6880 1550 6900 1650
rect 6830 1530 6900 1550
rect 7110 1650 7180 1670
rect 7110 1550 7130 1650
rect 7160 1550 7180 1650
rect 7220 1630 7240 1670
rect 7260 1630 7280 1670
rect 7220 1610 7280 1630
rect 7110 1530 7180 1550
rect 8170 1830 8250 1850
rect 7830 1800 7920 1820
rect 7830 1660 7850 1800
rect 7900 1660 7920 1800
rect 7830 1640 7920 1660
rect 8170 1630 8190 1830
rect 8230 1630 8250 1830
rect 8170 1610 8250 1630
rect 10740 1950 10800 1980
rect 10210 1670 10280 1690
rect 10210 1570 10230 1670
rect 10260 1570 10280 1670
rect 10210 1550 10280 1570
rect 10490 1670 10560 1690
rect 10490 1570 10510 1670
rect 10540 1570 10560 1670
rect 10490 1550 10560 1570
rect 10740 1530 10760 1950
rect 10780 1530 10800 1950
rect 10740 1500 10800 1530
rect 11250 1670 11320 1690
rect 11250 1570 11270 1670
rect 11300 1570 11320 1670
rect 11250 1550 11320 1570
rect 11530 1670 11600 1690
rect 11530 1570 11550 1670
rect 11580 1570 11600 1670
rect 11530 1550 11600 1570
rect 11810 1670 11880 1690
rect 11810 1570 11830 1670
rect 11860 1570 11880 1670
rect 11810 1550 11880 1570
rect 12100 1670 12170 1690
rect 12100 1570 12120 1670
rect 12150 1570 12170 1670
rect 12100 1550 12170 1570
<< nsubdiff >>
rect 2740 1930 2800 1960
rect 2210 1900 2280 1920
rect 2210 1800 2230 1900
rect 2260 1800 2280 1900
rect 2210 1780 2280 1800
rect 2490 1900 2560 1920
rect 2490 1800 2510 1900
rect 2540 1800 2560 1900
rect 2490 1780 2560 1800
rect 2740 1510 2760 1930
rect 2780 1510 2800 1930
rect 2740 1480 2800 1510
rect 3240 1900 3310 1920
rect 3240 1800 3260 1900
rect 3290 1800 3310 1900
rect 3240 1780 3310 1800
rect 3530 1900 3600 1920
rect 3530 1800 3550 1900
rect 3580 1800 3600 1900
rect 3530 1780 3600 1800
rect 3810 1900 3880 1920
rect 3810 1800 3830 1900
rect 3860 1800 3880 1900
rect 3810 1780 3880 1800
rect 4100 1900 4170 1920
rect 4100 1800 4120 1900
rect 4150 1800 4170 1900
rect 4100 1780 4170 1800
rect 5760 1930 5820 1960
rect 5230 1900 5300 1920
rect 5230 1800 5250 1900
rect 5280 1800 5300 1900
rect 5230 1780 5300 1800
rect 5510 1900 5580 1920
rect 5510 1800 5530 1900
rect 5560 1800 5580 1900
rect 5510 1780 5580 1800
rect 5760 1510 5780 1930
rect 5800 1510 5820 1930
rect 5760 1480 5820 1510
rect 6260 1900 6330 1920
rect 6260 1800 6280 1900
rect 6310 1800 6330 1900
rect 6260 1780 6330 1800
rect 6540 1900 6610 1920
rect 6540 1800 6560 1900
rect 6590 1800 6610 1900
rect 6540 1780 6610 1800
rect 6830 1900 6900 1920
rect 6830 1800 6850 1900
rect 6880 1800 6900 1900
rect 6830 1780 6900 1800
rect 7110 1900 7180 1920
rect 7110 1800 7130 1900
rect 7160 1800 7180 1900
rect 7500 1890 7560 1920
rect 7110 1780 7180 1800
rect 7500 1470 7520 1890
rect 7540 1470 7560 1890
rect 7500 1440 7560 1470
rect 8840 1900 8900 1930
rect 8530 1830 8610 1850
rect 8530 1630 8550 1830
rect 8590 1630 8610 1830
rect 8530 1610 8610 1630
rect 7940 1490 8000 1500
rect 7940 1470 7960 1490
rect 7980 1470 8000 1490
rect 7940 1460 8000 1470
rect 8840 1480 8860 1900
rect 8880 1480 8900 1900
rect 8840 1450 8900 1480
rect 10210 1920 10280 1940
rect 10210 1820 10230 1920
rect 10260 1820 10280 1920
rect 10210 1800 10280 1820
rect 10490 1920 10560 1940
rect 10490 1820 10510 1920
rect 10540 1820 10560 1920
rect 10490 1800 10560 1820
rect 11250 1920 11320 1940
rect 11250 1820 11270 1920
rect 11300 1820 11320 1920
rect 11250 1800 11320 1820
rect 11530 1920 11600 1940
rect 11530 1820 11550 1920
rect 11580 1820 11600 1920
rect 11530 1800 11600 1820
rect 11810 1920 11880 1940
rect 11810 1820 11830 1920
rect 11860 1820 11880 1920
rect 11810 1800 11880 1820
rect 12100 1920 12170 1940
rect 12100 1820 12120 1920
rect 12150 1820 12170 1920
rect 12100 1800 12170 1820
<< psubdiffcont >>
rect 2230 1550 2260 1650
rect 2510 1550 2540 1650
rect 3260 1550 3290 1650
rect 3550 1550 3580 1650
rect 3830 1550 3860 1650
rect 4120 1550 4150 1650
rect 5250 1550 5280 1650
rect 5530 1550 5560 1650
rect 7240 1770 7260 1810
rect 6280 1550 6310 1650
rect 6560 1550 6590 1650
rect 6850 1550 6880 1650
rect 7130 1550 7160 1650
rect 7240 1630 7260 1670
rect 7850 1660 7900 1800
rect 8190 1630 8230 1830
rect 10230 1570 10260 1670
rect 10510 1570 10540 1670
rect 10760 1530 10780 1950
rect 11270 1570 11300 1670
rect 11550 1570 11580 1670
rect 11830 1570 11860 1670
rect 12120 1570 12150 1670
<< nsubdiffcont >>
rect 2230 1800 2260 1900
rect 2510 1800 2540 1900
rect 2760 1510 2780 1930
rect 3260 1800 3290 1900
rect 3550 1800 3580 1900
rect 3830 1800 3860 1900
rect 4120 1800 4150 1900
rect 5250 1800 5280 1900
rect 5530 1800 5560 1900
rect 5780 1510 5800 1930
rect 6280 1800 6310 1900
rect 6560 1800 6590 1900
rect 6850 1800 6880 1900
rect 7130 1800 7160 1900
rect 7520 1470 7540 1890
rect 8550 1630 8590 1830
rect 7960 1470 7980 1490
rect 8860 1480 8880 1900
rect 10230 1820 10260 1920
rect 10510 1820 10540 1920
rect 11270 1820 11300 1920
rect 11550 1820 11580 1920
rect 11830 1820 11860 1920
rect 12120 1820 12150 1920
<< poly >>
rect 5900 2000 5940 2010
rect 1160 1980 2920 2000
rect 1160 1500 1210 1980
rect 1910 1500 1960 1980
rect 2880 1960 2920 1980
rect 4220 1980 5940 2000
rect 2100 1920 2140 1950
rect 2380 1920 2420 1950
rect 2100 1760 2140 1780
rect 2380 1760 2420 1780
rect 2100 1670 2140 1690
rect 2380 1670 2420 1690
rect 2100 1490 2140 1530
rect 2380 1490 2420 1530
rect 3130 1920 3170 1960
rect 3420 1920 3460 1960
rect 3700 1920 3740 1960
rect 3990 1920 4030 1960
rect 3130 1760 3170 1780
rect 3420 1760 3460 1780
rect 3700 1760 3740 1780
rect 3990 1760 4030 1780
rect 3130 1670 3170 1690
rect 3420 1670 3460 1690
rect 3700 1670 3740 1690
rect 3990 1670 4030 1690
rect 3130 1490 3170 1530
rect 3420 1490 3460 1530
rect 3700 1490 3740 1530
rect 3990 1490 4030 1530
rect 4220 1500 4270 1980
rect 4970 1500 5020 1980
rect 5900 1960 5940 1980
rect 9160 2000 10920 2020
rect 5120 1920 5160 1950
rect 5400 1920 5440 1950
rect 5120 1760 5160 1780
rect 5400 1760 5440 1780
rect 5120 1670 5160 1690
rect 5400 1670 5440 1690
rect 2880 1470 2920 1480
rect 2560 1450 2590 1470
rect 2680 1450 2920 1470
rect 2880 1430 2920 1450
rect 5120 1490 5160 1530
rect 5400 1490 5440 1530
rect 6150 1920 6190 1960
rect 6430 1920 6470 1960
rect 6720 1920 6760 1960
rect 7000 1920 7040 1960
rect 7640 1920 7680 1970
rect 8980 1930 9020 1970
rect 7330 1830 7370 1850
rect 6150 1760 6190 1780
rect 6430 1760 6470 1780
rect 6720 1760 6760 1780
rect 7000 1760 7040 1780
rect 7330 1730 7370 1750
rect 7330 1710 7340 1730
rect 7360 1710 7370 1730
rect 7330 1690 7370 1710
rect 6150 1670 6190 1690
rect 6430 1670 6470 1690
rect 6720 1670 6760 1690
rect 7000 1670 7040 1690
rect 7330 1570 7370 1610
rect 6150 1490 6190 1530
rect 6430 1490 6470 1530
rect 6720 1490 6760 1530
rect 7000 1490 7040 1530
rect 5900 1470 5940 1480
rect 5580 1450 5610 1470
rect 5700 1450 5940 1470
rect 5900 1430 5940 1450
rect 8330 1900 8370 1910
rect 8330 1880 8340 1900
rect 8360 1880 8370 1900
rect 8010 1820 8050 1870
rect 8330 1850 8370 1880
rect 8690 1900 8730 1910
rect 8690 1880 8700 1900
rect 8720 1880 8730 1900
rect 8690 1850 8730 1880
rect 8010 1620 8050 1640
rect 8010 1600 8020 1620
rect 8040 1600 8050 1620
rect 8010 1590 8050 1600
rect 8330 1580 8370 1610
rect 8690 1580 8730 1610
rect 8060 1500 8100 1540
rect 8060 1440 8100 1460
rect 9160 1520 9210 2000
rect 9910 1520 9960 2000
rect 10880 1980 10920 2000
rect 10100 1940 10140 1970
rect 10380 1940 10420 1970
rect 10100 1780 10140 1800
rect 10380 1780 10420 1800
rect 10100 1690 10140 1710
rect 10380 1690 10420 1710
rect 10100 1510 10140 1550
rect 10380 1510 10420 1550
rect 11140 1940 11180 1980
rect 11420 1940 11460 1980
rect 11700 1940 11740 1980
rect 11990 1940 12030 1980
rect 11140 1780 11180 1800
rect 11420 1780 11460 1800
rect 11700 1780 11740 1800
rect 11990 1780 12030 1800
rect 11140 1690 11180 1710
rect 11420 1690 11460 1710
rect 11700 1690 11740 1710
rect 11990 1690 12030 1710
rect 11140 1510 11180 1550
rect 11420 1510 11460 1550
rect 11700 1510 11740 1550
rect 11990 1510 12030 1550
rect 10880 1490 10920 1500
rect 10580 1470 10610 1490
rect 10700 1470 10920 1490
rect 7640 1430 7680 1440
rect 8000 1430 8100 1440
rect 8980 1430 9020 1450
rect 7640 1410 8020 1430
rect 8040 1410 9020 1430
rect 10880 1450 10920 1470
rect 8000 1400 8060 1410
<< polycont >>
rect 7340 1710 7360 1730
rect 8340 1880 8360 1900
rect 8700 1880 8720 1900
rect 8020 1600 8040 1620
rect 8020 1410 8040 1430
<< locali >>
rect 10750 1950 10790 1970
rect 2750 1930 2790 1950
rect 2040 1900 2090 1910
rect 2040 1800 2050 1900
rect 2080 1800 2090 1900
rect 2040 1790 2090 1800
rect 2150 1900 2200 1910
rect 2150 1800 2160 1900
rect 2190 1800 2200 1900
rect 2150 1790 2200 1800
rect 2220 1900 2270 1910
rect 2220 1800 2230 1900
rect 2260 1800 2270 1900
rect 2220 1790 2270 1800
rect 2320 1900 2370 1910
rect 2320 1800 2330 1900
rect 2360 1800 2370 1900
rect 2320 1790 2370 1800
rect 2430 1900 2480 1910
rect 2430 1800 2440 1900
rect 2470 1800 2480 1900
rect 2430 1790 2480 1800
rect 2500 1900 2550 1910
rect 2500 1800 2510 1900
rect 2540 1800 2550 1900
rect 2500 1790 2550 1800
rect 2040 1650 2090 1660
rect 2040 1550 2050 1650
rect 2080 1550 2090 1650
rect 2040 1540 2090 1550
rect 2150 1650 2200 1660
rect 2150 1550 2160 1650
rect 2190 1550 2200 1650
rect 2150 1540 2200 1550
rect 2220 1650 2270 1660
rect 2220 1550 2230 1650
rect 2260 1550 2270 1650
rect 2220 1540 2270 1550
rect 2320 1650 2370 1660
rect 2320 1550 2330 1650
rect 2360 1550 2370 1650
rect 2320 1540 2370 1550
rect 2430 1650 2480 1660
rect 2430 1550 2440 1650
rect 2470 1550 2480 1650
rect 2430 1540 2480 1550
rect 2500 1650 2550 1660
rect 2500 1550 2510 1650
rect 2540 1550 2550 1650
rect 2500 1540 2550 1550
rect 2750 1510 2760 1930
rect 2780 1510 2790 1930
rect 2750 1490 2790 1510
rect 2820 1930 2860 1950
rect 2820 1510 2830 1930
rect 2850 1510 2860 1930
rect 2820 1490 2860 1510
rect 2940 1930 2980 1950
rect 2940 1510 2950 1930
rect 2970 1510 2980 1930
rect 5770 1930 5810 1950
rect 3070 1900 3120 1910
rect 3070 1800 3080 1900
rect 3110 1800 3120 1900
rect 3070 1790 3120 1800
rect 3180 1900 3230 1910
rect 3180 1800 3190 1900
rect 3220 1800 3230 1900
rect 3180 1790 3230 1800
rect 3250 1900 3300 1910
rect 3250 1800 3260 1900
rect 3290 1800 3300 1900
rect 3250 1790 3300 1800
rect 3360 1900 3410 1910
rect 3360 1800 3370 1900
rect 3400 1800 3410 1900
rect 3360 1790 3410 1800
rect 3470 1900 3520 1910
rect 3470 1800 3480 1900
rect 3510 1800 3520 1900
rect 3470 1790 3520 1800
rect 3540 1900 3590 1910
rect 3540 1800 3550 1900
rect 3580 1800 3590 1900
rect 3540 1790 3590 1800
rect 3640 1900 3690 1910
rect 3640 1800 3650 1900
rect 3680 1800 3690 1900
rect 3640 1790 3690 1800
rect 3750 1900 3800 1910
rect 3750 1800 3760 1900
rect 3790 1800 3800 1900
rect 3750 1790 3800 1800
rect 3820 1900 3870 1910
rect 3820 1800 3830 1900
rect 3860 1800 3870 1900
rect 3820 1790 3870 1800
rect 3930 1900 3980 1910
rect 3930 1800 3940 1900
rect 3970 1800 3980 1900
rect 3930 1790 3980 1800
rect 4040 1900 4090 1910
rect 4040 1800 4050 1900
rect 4080 1800 4090 1900
rect 4040 1790 4090 1800
rect 4110 1900 4160 1910
rect 4110 1800 4120 1900
rect 4150 1800 4160 1900
rect 4110 1790 4160 1800
rect 5060 1900 5110 1910
rect 5060 1800 5070 1900
rect 5100 1800 5110 1900
rect 5060 1790 5110 1800
rect 5170 1900 5220 1910
rect 5170 1800 5180 1900
rect 5210 1800 5220 1900
rect 5170 1790 5220 1800
rect 5240 1900 5290 1910
rect 5240 1800 5250 1900
rect 5280 1800 5290 1900
rect 5240 1790 5290 1800
rect 5340 1900 5390 1910
rect 5340 1800 5350 1900
rect 5380 1800 5390 1900
rect 5340 1790 5390 1800
rect 5450 1900 5500 1910
rect 5450 1800 5460 1900
rect 5490 1800 5500 1900
rect 5450 1790 5500 1800
rect 5520 1900 5570 1910
rect 5520 1800 5530 1900
rect 5560 1800 5570 1900
rect 5520 1790 5570 1800
rect 3070 1650 3120 1660
rect 3070 1550 3080 1650
rect 3110 1550 3120 1650
rect 3070 1540 3120 1550
rect 3180 1650 3230 1660
rect 3180 1550 3190 1650
rect 3220 1550 3230 1650
rect 3180 1540 3230 1550
rect 3250 1650 3300 1660
rect 3250 1550 3260 1650
rect 3290 1550 3300 1650
rect 3250 1540 3300 1550
rect 3360 1650 3410 1660
rect 3360 1550 3370 1650
rect 3400 1550 3410 1650
rect 3360 1540 3410 1550
rect 3470 1650 3520 1660
rect 3470 1550 3480 1650
rect 3510 1550 3520 1650
rect 3470 1540 3520 1550
rect 3540 1650 3590 1660
rect 3540 1550 3550 1650
rect 3580 1550 3590 1650
rect 3540 1540 3590 1550
rect 3640 1650 3690 1660
rect 3640 1550 3650 1650
rect 3680 1550 3690 1650
rect 3640 1540 3690 1550
rect 3750 1650 3800 1660
rect 3750 1550 3760 1650
rect 3790 1550 3800 1650
rect 3750 1540 3800 1550
rect 3820 1650 3870 1660
rect 3820 1550 3830 1650
rect 3860 1550 3870 1650
rect 3820 1540 3870 1550
rect 3930 1650 3980 1660
rect 3930 1550 3940 1650
rect 3970 1550 3980 1650
rect 3930 1540 3980 1550
rect 4040 1650 4090 1660
rect 4040 1550 4050 1650
rect 4080 1550 4090 1650
rect 4040 1540 4090 1550
rect 4110 1650 4160 1660
rect 4110 1550 4120 1650
rect 4150 1550 4160 1650
rect 4110 1540 4160 1550
rect 5060 1650 5110 1660
rect 5060 1550 5070 1650
rect 5100 1550 5110 1650
rect 5060 1540 5110 1550
rect 5170 1650 5220 1660
rect 5170 1550 5180 1650
rect 5210 1550 5220 1650
rect 5170 1540 5220 1550
rect 5240 1650 5290 1660
rect 5240 1550 5250 1650
rect 5280 1550 5290 1650
rect 5240 1540 5290 1550
rect 5340 1650 5390 1660
rect 5340 1550 5350 1650
rect 5380 1550 5390 1650
rect 5340 1540 5390 1550
rect 5450 1650 5500 1660
rect 5450 1550 5460 1650
rect 5490 1550 5500 1650
rect 5450 1540 5500 1550
rect 5520 1650 5570 1660
rect 5520 1550 5530 1650
rect 5560 1550 5570 1650
rect 5520 1540 5570 1550
rect 2940 1490 2980 1510
rect 5770 1510 5780 1930
rect 5800 1510 5810 1930
rect 5770 1490 5810 1510
rect 5840 1930 5880 1950
rect 5840 1510 5850 1930
rect 5870 1510 5880 1930
rect 5840 1490 5880 1510
rect 5960 1930 6000 1950
rect 5960 1510 5970 1930
rect 5990 1510 6000 1930
rect 10040 1920 10090 1930
rect 6090 1900 6140 1910
rect 6090 1800 6100 1900
rect 6130 1800 6140 1900
rect 6090 1790 6140 1800
rect 6200 1900 6250 1910
rect 6200 1800 6210 1900
rect 6240 1800 6250 1900
rect 6200 1790 6250 1800
rect 6270 1900 6320 1910
rect 6270 1800 6280 1900
rect 6310 1800 6320 1900
rect 6270 1790 6320 1800
rect 6370 1900 6420 1910
rect 6370 1800 6380 1900
rect 6410 1800 6420 1900
rect 6370 1790 6420 1800
rect 6480 1900 6530 1910
rect 6480 1800 6490 1900
rect 6520 1800 6530 1900
rect 6480 1790 6530 1800
rect 6550 1900 6600 1910
rect 6550 1800 6560 1900
rect 6590 1800 6600 1900
rect 6550 1790 6600 1800
rect 6660 1900 6710 1910
rect 6660 1800 6670 1900
rect 6700 1800 6710 1900
rect 6660 1790 6710 1800
rect 6770 1900 6820 1910
rect 6770 1800 6780 1900
rect 6810 1800 6820 1900
rect 6770 1790 6820 1800
rect 6840 1900 6890 1910
rect 6840 1800 6850 1900
rect 6880 1800 6890 1900
rect 6840 1790 6890 1800
rect 6940 1900 6990 1910
rect 6940 1800 6950 1900
rect 6980 1800 6990 1900
rect 6940 1790 6990 1800
rect 7050 1900 7100 1910
rect 7050 1800 7060 1900
rect 7090 1800 7100 1900
rect 7050 1790 7100 1800
rect 7120 1900 7170 1910
rect 7120 1800 7130 1900
rect 7160 1800 7170 1900
rect 7510 1890 7550 1910
rect 7120 1790 7170 1800
rect 7230 1810 7270 1820
rect 7230 1770 7240 1810
rect 7260 1770 7270 1810
rect 7230 1760 7270 1770
rect 7290 1810 7320 1820
rect 7290 1770 7300 1810
rect 7290 1760 7320 1770
rect 7380 1810 7420 1820
rect 7380 1770 7390 1810
rect 7410 1770 7420 1810
rect 7380 1760 7420 1770
rect 7330 1730 7370 1740
rect 7330 1710 7340 1730
rect 7360 1710 7370 1730
rect 7330 1700 7370 1710
rect 7230 1670 7270 1680
rect 6090 1650 6140 1660
rect 6090 1550 6100 1650
rect 6130 1550 6140 1650
rect 6090 1540 6140 1550
rect 6200 1650 6250 1660
rect 6200 1550 6210 1650
rect 6240 1550 6250 1650
rect 6200 1540 6250 1550
rect 6270 1650 6320 1660
rect 6270 1550 6280 1650
rect 6310 1550 6320 1650
rect 6270 1540 6320 1550
rect 6370 1650 6420 1660
rect 6370 1550 6380 1650
rect 6410 1550 6420 1650
rect 6370 1540 6420 1550
rect 6480 1650 6530 1660
rect 6480 1550 6490 1650
rect 6520 1550 6530 1650
rect 6480 1540 6530 1550
rect 6550 1650 6600 1660
rect 6550 1550 6560 1650
rect 6590 1550 6600 1650
rect 6550 1540 6600 1550
rect 6660 1650 6710 1660
rect 6660 1550 6670 1650
rect 6700 1550 6710 1650
rect 6660 1540 6710 1550
rect 6770 1650 6820 1660
rect 6770 1550 6780 1650
rect 6810 1550 6820 1650
rect 6770 1540 6820 1550
rect 6840 1650 6890 1660
rect 6840 1550 6850 1650
rect 6880 1550 6890 1650
rect 6840 1540 6890 1550
rect 6940 1650 6990 1660
rect 6940 1550 6950 1650
rect 6980 1550 6990 1650
rect 6940 1540 6990 1550
rect 7050 1650 7100 1660
rect 7050 1550 7060 1650
rect 7090 1550 7100 1650
rect 7050 1540 7100 1550
rect 7120 1650 7170 1660
rect 7120 1550 7130 1650
rect 7160 1550 7170 1650
rect 7230 1630 7240 1670
rect 7260 1630 7270 1670
rect 7230 1620 7270 1630
rect 7290 1670 7320 1680
rect 7290 1630 7300 1670
rect 7290 1620 7320 1630
rect 7380 1670 7420 1680
rect 7380 1630 7390 1670
rect 7410 1630 7420 1670
rect 7380 1620 7420 1630
rect 7120 1540 7170 1550
rect 5960 1490 6000 1510
rect 1230 1470 1890 1480
rect 1230 1430 1670 1470
rect 1730 1430 1810 1470
rect 1870 1430 1890 1470
rect 4290 1470 4950 1480
rect 4290 1440 4730 1470
rect 4790 1440 4870 1470
rect 4930 1440 4950 1470
rect 7510 1470 7520 1890
rect 7540 1470 7550 1890
rect 7510 1450 7550 1470
rect 7580 1890 7620 1910
rect 7580 1470 7590 1890
rect 7610 1470 7620 1890
rect 7580 1450 7620 1470
rect 7700 1890 7740 1910
rect 7700 1470 7710 1890
rect 7730 1470 7740 1890
rect 8330 1900 8370 1910
rect 8330 1880 8340 1900
rect 8360 1880 8370 1900
rect 8330 1860 8370 1880
rect 8690 1900 8730 1910
rect 8690 1880 8700 1900
rect 8720 1880 8730 1900
rect 8690 1860 8730 1880
rect 8850 1900 8890 1920
rect 8180 1830 8240 1840
rect 7840 1800 7910 1810
rect 7840 1660 7850 1800
rect 7900 1660 7910 1800
rect 7840 1650 7910 1660
rect 7930 1800 8000 1810
rect 7930 1660 7940 1800
rect 7990 1660 8000 1800
rect 7930 1650 8000 1660
rect 8060 1800 8130 1810
rect 8060 1660 8070 1800
rect 8120 1660 8130 1800
rect 8060 1650 8130 1660
rect 8180 1630 8190 1830
rect 8230 1630 8240 1830
rect 8010 1620 8050 1630
rect 8180 1620 8240 1630
rect 8260 1830 8320 1840
rect 8260 1630 8270 1830
rect 8310 1630 8320 1830
rect 8260 1620 8320 1630
rect 8380 1830 8440 1840
rect 8380 1630 8390 1830
rect 8430 1630 8440 1830
rect 8380 1620 8440 1630
rect 8540 1830 8600 1840
rect 8540 1630 8550 1830
rect 8590 1630 8600 1830
rect 8540 1620 8600 1630
rect 8620 1830 8680 1840
rect 8620 1630 8630 1830
rect 8670 1630 8680 1830
rect 8620 1620 8680 1630
rect 8740 1830 8800 1840
rect 8740 1630 8750 1830
rect 8790 1630 8800 1830
rect 8740 1620 8800 1630
rect 8010 1600 8020 1620
rect 8040 1600 8050 1620
rect 8010 1590 8050 1600
rect 7950 1470 7960 1490
rect 7980 1470 7990 1490
rect 8010 1470 8020 1490
rect 8040 1470 8050 1490
rect 8110 1470 8120 1490
rect 8140 1470 8150 1490
rect 8850 1480 8860 1900
rect 8880 1480 8890 1900
rect 7700 1450 7740 1470
rect 8850 1460 8890 1480
rect 8920 1900 8960 1920
rect 8920 1480 8930 1900
rect 8950 1480 8960 1900
rect 8920 1460 8960 1480
rect 9040 1900 9080 1920
rect 9040 1480 9050 1900
rect 9070 1480 9080 1900
rect 10040 1820 10050 1920
rect 10080 1820 10090 1920
rect 10040 1810 10090 1820
rect 10150 1920 10200 1930
rect 10150 1820 10160 1920
rect 10190 1820 10200 1920
rect 10150 1810 10200 1820
rect 10220 1920 10270 1930
rect 10220 1820 10230 1920
rect 10260 1820 10270 1920
rect 10220 1810 10270 1820
rect 10320 1920 10370 1930
rect 10320 1820 10330 1920
rect 10360 1820 10370 1920
rect 10320 1810 10370 1820
rect 10430 1920 10480 1930
rect 10430 1820 10440 1920
rect 10470 1820 10480 1920
rect 10430 1810 10480 1820
rect 10500 1920 10550 1930
rect 10500 1820 10510 1920
rect 10540 1820 10550 1920
rect 10500 1810 10550 1820
rect 10040 1670 10090 1680
rect 10040 1570 10050 1670
rect 10080 1570 10090 1670
rect 10040 1560 10090 1570
rect 10150 1670 10200 1680
rect 10150 1570 10160 1670
rect 10190 1570 10200 1670
rect 10150 1560 10200 1570
rect 10220 1670 10270 1680
rect 10220 1570 10230 1670
rect 10260 1570 10270 1670
rect 10220 1560 10270 1570
rect 10320 1670 10370 1680
rect 10320 1570 10330 1670
rect 10360 1570 10370 1670
rect 10320 1560 10370 1570
rect 10430 1670 10480 1680
rect 10430 1570 10440 1670
rect 10470 1570 10480 1670
rect 10430 1560 10480 1570
rect 10500 1670 10550 1680
rect 10500 1570 10510 1670
rect 10540 1570 10550 1670
rect 10500 1560 10550 1570
rect 10750 1530 10760 1950
rect 10780 1530 10790 1950
rect 10750 1510 10790 1530
rect 10820 1950 10860 1970
rect 10820 1530 10830 1950
rect 10850 1530 10860 1950
rect 10820 1510 10860 1530
rect 10940 1950 10980 1970
rect 10940 1530 10950 1950
rect 10970 1530 10980 1950
rect 11080 1920 11130 1930
rect 11080 1820 11090 1920
rect 11120 1820 11130 1920
rect 11080 1810 11130 1820
rect 11190 1920 11240 1930
rect 11190 1820 11200 1920
rect 11230 1820 11240 1920
rect 11190 1810 11240 1820
rect 11260 1920 11310 1930
rect 11260 1820 11270 1920
rect 11300 1820 11310 1920
rect 11260 1810 11310 1820
rect 11360 1920 11410 1930
rect 11360 1820 11370 1920
rect 11400 1820 11410 1920
rect 11360 1810 11410 1820
rect 11470 1920 11520 1930
rect 11470 1820 11480 1920
rect 11510 1820 11520 1920
rect 11470 1810 11520 1820
rect 11540 1920 11590 1930
rect 11540 1820 11550 1920
rect 11580 1820 11590 1920
rect 11540 1810 11590 1820
rect 11640 1920 11690 1930
rect 11640 1820 11650 1920
rect 11680 1820 11690 1920
rect 11640 1810 11690 1820
rect 11750 1920 11800 1930
rect 11750 1820 11760 1920
rect 11790 1820 11800 1920
rect 11750 1810 11800 1820
rect 11820 1920 11870 1930
rect 11820 1820 11830 1920
rect 11860 1820 11870 1920
rect 11820 1810 11870 1820
rect 11930 1920 11980 1930
rect 11930 1820 11940 1920
rect 11970 1820 11980 1920
rect 11930 1810 11980 1820
rect 12040 1920 12090 1930
rect 12040 1820 12050 1920
rect 12080 1820 12090 1920
rect 12040 1810 12090 1820
rect 12110 1920 12160 1930
rect 12110 1820 12120 1920
rect 12150 1820 12160 1920
rect 12110 1810 12160 1820
rect 11080 1670 11130 1680
rect 11080 1570 11090 1670
rect 11120 1570 11130 1670
rect 11080 1560 11130 1570
rect 11190 1670 11240 1680
rect 11190 1570 11200 1670
rect 11230 1570 11240 1670
rect 11190 1560 11240 1570
rect 11260 1670 11310 1680
rect 11260 1570 11270 1670
rect 11300 1570 11310 1670
rect 11260 1560 11310 1570
rect 11360 1670 11410 1680
rect 11360 1570 11370 1670
rect 11400 1570 11410 1670
rect 11360 1560 11410 1570
rect 11470 1670 11520 1680
rect 11470 1570 11480 1670
rect 11510 1570 11520 1670
rect 11470 1560 11520 1570
rect 11540 1670 11590 1680
rect 11540 1570 11550 1670
rect 11580 1570 11590 1670
rect 11540 1560 11590 1570
rect 11640 1670 11690 1680
rect 11640 1570 11650 1670
rect 11680 1570 11690 1670
rect 11640 1560 11690 1570
rect 11750 1670 11800 1680
rect 11750 1570 11760 1670
rect 11790 1570 11800 1670
rect 11750 1560 11800 1570
rect 11820 1670 11870 1680
rect 11820 1570 11830 1670
rect 11860 1570 11870 1670
rect 11820 1560 11870 1570
rect 11930 1670 11980 1680
rect 11930 1570 11940 1670
rect 11970 1570 11980 1670
rect 11930 1560 11980 1570
rect 12040 1670 12090 1680
rect 12040 1570 12050 1670
rect 12080 1570 12090 1670
rect 12040 1560 12090 1570
rect 12110 1670 12160 1680
rect 12110 1570 12120 1670
rect 12150 1570 12160 1670
rect 12110 1560 12160 1570
rect 10940 1510 10980 1530
rect 9040 1460 9080 1480
rect 9230 1490 9890 1500
rect 9230 1450 9670 1490
rect 9730 1450 9810 1490
rect 9870 1450 9890 1490
rect 9230 1440 9890 1450
rect 4290 1430 4950 1440
rect 8010 1430 8050 1440
rect 1230 1420 1890 1430
rect 8010 1410 8020 1430
rect 8040 1410 8050 1430
rect 8010 1400 8050 1410
<< viali >>
rect 2050 1840 2080 1860
rect 2160 1840 2190 1860
rect 2230 1860 2260 1880
rect 2330 1840 2360 1860
rect 2440 1840 2470 1860
rect 2510 1850 2540 1870
rect 2050 1580 2080 1600
rect 2160 1580 2190 1600
rect 2230 1580 2260 1600
rect 2330 1580 2360 1600
rect 2440 1580 2470 1600
rect 2510 1570 2540 1590
rect 2610 1580 2620 1600
rect 2620 1580 2640 1600
rect 2640 1580 2650 1600
rect 2610 1570 2650 1580
rect 2760 1880 2780 1900
rect 2830 1700 2850 1720
rect 2950 1520 2970 1540
rect 3080 1840 3110 1860
rect 3190 1840 3220 1860
rect 3260 1840 3290 1860
rect 3370 1840 3400 1860
rect 3480 1840 3510 1860
rect 3550 1840 3580 1860
rect 3650 1840 3680 1860
rect 3760 1840 3790 1860
rect 3830 1840 3860 1860
rect 3940 1840 3970 1860
rect 4050 1840 4080 1860
rect 4120 1840 4150 1860
rect 5070 1840 5100 1860
rect 5180 1840 5210 1860
rect 5250 1840 5280 1860
rect 5350 1840 5380 1860
rect 5460 1840 5490 1860
rect 5530 1850 5560 1870
rect 3080 1580 3110 1600
rect 3190 1580 3220 1600
rect 3260 1570 3290 1590
rect 3370 1580 3400 1600
rect 3480 1580 3510 1600
rect 3550 1570 3580 1590
rect 3650 1580 3680 1600
rect 3760 1580 3790 1600
rect 3830 1570 3860 1590
rect 3940 1580 3970 1600
rect 4050 1580 4080 1600
rect 4120 1570 4150 1590
rect 5070 1580 5100 1600
rect 5180 1580 5210 1600
rect 5250 1570 5280 1590
rect 5350 1580 5380 1600
rect 5460 1580 5490 1600
rect 5530 1570 5560 1590
rect 5640 1580 5650 1600
rect 5650 1580 5670 1600
rect 5670 1580 5680 1600
rect 5640 1570 5680 1580
rect 5780 1840 5800 1860
rect 5850 1700 5870 1720
rect 5970 1520 5990 1540
rect 6100 1840 6130 1860
rect 6210 1840 6240 1860
rect 6280 1850 6310 1870
rect 6380 1840 6410 1860
rect 6490 1840 6520 1860
rect 6560 1850 6590 1870
rect 6670 1840 6700 1860
rect 6780 1840 6810 1860
rect 6850 1840 6880 1860
rect 6950 1840 6980 1860
rect 7060 1840 7090 1860
rect 7130 1840 7160 1860
rect 7240 1770 7260 1810
rect 7300 1771 7317 1791
rect 7390 1770 7410 1810
rect 7340 1710 7360 1730
rect 6100 1580 6130 1600
rect 6210 1580 6240 1600
rect 6280 1570 6310 1590
rect 6380 1580 6410 1600
rect 6490 1580 6520 1600
rect 6560 1570 6590 1590
rect 6670 1580 6700 1600
rect 6780 1580 6810 1600
rect 6850 1570 6880 1590
rect 6950 1580 6980 1600
rect 7060 1580 7090 1600
rect 7130 1570 7160 1590
rect 7240 1630 7260 1650
rect 7300 1630 7317 1650
rect 7390 1630 7410 1670
rect 1670 1430 1730 1470
rect 1810 1430 1870 1470
rect 4730 1440 4790 1470
rect 4870 1440 4930 1470
rect 7520 1750 7540 1770
rect 7590 1770 7610 1790
rect 7710 1850 7730 1880
rect 8340 1880 8360 1900
rect 8700 1880 8720 1900
rect 7860 1680 7890 1700
rect 7950 1690 7980 1720
rect 8080 1770 8110 1800
rect 8190 1660 8230 1680
rect 8270 1670 8310 1700
rect 8390 1780 8430 1810
rect 8550 1690 8590 1720
rect 8630 1780 8670 1810
rect 8750 1710 8790 1740
rect 8020 1600 8040 1620
rect 8020 1490 8040 1492
rect 7960 1470 7980 1490
rect 8020 1474 8040 1490
rect 8120 1470 8140 1490
rect 8860 1840 8880 1860
rect 9050 1830 9070 1860
rect 10050 1860 10080 1880
rect 10160 1860 10190 1880
rect 10230 1870 10260 1890
rect 10330 1860 10360 1880
rect 10440 1860 10470 1880
rect 10510 1870 10540 1890
rect 10050 1600 10080 1620
rect 10160 1600 10190 1620
rect 10230 1590 10260 1610
rect 10330 1600 10360 1620
rect 10440 1600 10470 1620
rect 10510 1590 10540 1610
rect 10640 1590 10650 1610
rect 10650 1590 10670 1610
rect 10670 1590 10680 1610
rect 10640 1580 10680 1590
rect 10760 1560 10780 1580
rect 10830 1720 10850 1740
rect 10950 1530 10970 1560
rect 11090 1860 11120 1880
rect 11200 1860 11230 1880
rect 11270 1870 11300 1890
rect 11370 1860 11400 1880
rect 11480 1860 11510 1880
rect 11550 1870 11580 1890
rect 11650 1860 11680 1880
rect 11760 1860 11790 1880
rect 11830 1860 11860 1880
rect 11940 1860 11970 1880
rect 12050 1860 12080 1880
rect 12120 1860 12150 1880
rect 11090 1600 11120 1620
rect 11200 1600 11230 1620
rect 11270 1590 11300 1610
rect 11370 1600 11400 1620
rect 11480 1600 11510 1620
rect 11550 1590 11580 1610
rect 11650 1600 11680 1620
rect 11760 1600 11790 1620
rect 11830 1590 11860 1610
rect 11940 1600 11970 1620
rect 12050 1600 12080 1620
rect 12120 1590 12150 1610
rect 9670 1450 9730 1490
rect 9810 1450 9870 1490
rect 8020 1410 8040 1430
<< metal1 >>
rect 3180 1990 7420 2010
rect 2040 1860 2090 1880
rect 2040 1840 2050 1860
rect 2080 1840 2090 1860
rect 2040 1600 2090 1840
rect 2040 1580 2050 1600
rect 2080 1580 2090 1600
rect 2040 1480 2090 1580
rect 2150 1860 2200 1970
rect 2150 1840 2160 1860
rect 2190 1840 2200 1860
rect 2150 1600 2200 1840
rect 2220 1880 2270 1910
rect 2220 1850 2230 1880
rect 2260 1850 2270 1880
rect 2220 1790 2270 1850
rect 2320 1860 2370 1880
rect 2320 1840 2330 1860
rect 2360 1840 2370 1860
rect 2150 1580 2160 1600
rect 2190 1580 2200 1600
rect 2150 1540 2200 1580
rect 2220 1610 2270 1660
rect 2220 1580 2230 1610
rect 2260 1580 2270 1610
rect 2220 1540 2270 1580
rect 2320 1600 2370 1840
rect 2320 1580 2330 1600
rect 2360 1580 2370 1600
rect 2320 1480 2370 1580
rect 2430 1860 2480 1970
rect 2430 1840 2440 1860
rect 2470 1840 2480 1860
rect 2430 1600 2480 1840
rect 2500 1870 2550 1910
rect 2500 1840 2510 1870
rect 2540 1840 2550 1870
rect 2500 1790 2550 1840
rect 2750 1901 2790 1950
rect 2750 1873 2754 1901
rect 2787 1873 2790 1901
rect 2750 1830 2790 1873
rect 3070 1860 3120 1910
rect 3070 1840 3080 1860
rect 3110 1840 3120 1860
rect 3070 1730 3120 1840
rect 2820 1720 3120 1730
rect 2820 1700 2830 1720
rect 2850 1700 3120 1720
rect 2820 1690 3120 1700
rect 2430 1580 2440 1600
rect 2470 1580 2480 1600
rect 2430 1540 2480 1580
rect 2500 1600 2550 1660
rect 2500 1570 2510 1600
rect 2540 1570 2550 1600
rect 2500 1540 2550 1570
rect 2600 1600 2660 1660
rect 2600 1560 2610 1600
rect 2650 1560 2660 1600
rect 2600 1540 2660 1560
rect 3070 1600 3120 1690
rect 3070 1580 3080 1600
rect 3110 1580 3120 1600
rect 2940 1540 2980 1550
rect 1640 1470 2370 1480
rect 1640 1430 1670 1470
rect 1730 1430 1810 1470
rect 1870 1430 2370 1470
rect 1640 1420 2370 1430
rect 2940 1520 2950 1540
rect 2970 1520 2980 1540
rect 2940 1410 2980 1520
rect 3070 1470 3120 1580
rect 3180 1860 3230 1990
rect 3180 1840 3190 1860
rect 3220 1840 3230 1860
rect 3180 1600 3230 1840
rect 3250 1860 3300 1910
rect 3250 1830 3260 1860
rect 3290 1830 3300 1860
rect 3250 1790 3300 1830
rect 3360 1860 3410 1880
rect 3360 1840 3370 1860
rect 3400 1840 3410 1860
rect 3180 1580 3190 1600
rect 3220 1580 3230 1600
rect 3180 1540 3230 1580
rect 3250 1600 3300 1660
rect 3250 1570 3260 1600
rect 3290 1570 3300 1600
rect 3250 1540 3300 1570
rect 3360 1600 3410 1840
rect 3360 1580 3370 1600
rect 3400 1580 3410 1600
rect 3360 1470 3410 1580
rect 3470 1860 3520 1910
rect 3470 1840 3480 1860
rect 3510 1840 3520 1860
rect 3470 1730 3520 1840
rect 3540 1860 3590 1910
rect 3540 1830 3550 1860
rect 3580 1830 3590 1860
rect 3540 1790 3590 1830
rect 3640 1860 3690 1880
rect 3640 1840 3650 1860
rect 3680 1840 3690 1860
rect 3640 1730 3690 1840
rect 3470 1690 3690 1730
rect 3470 1600 3520 1690
rect 3470 1580 3480 1600
rect 3510 1580 3520 1600
rect 3470 1540 3520 1580
rect 3540 1600 3590 1660
rect 3540 1570 3550 1600
rect 3580 1570 3590 1600
rect 3540 1540 3590 1570
rect 3640 1600 3690 1690
rect 3640 1580 3650 1600
rect 3680 1580 3690 1600
rect 3070 1450 3410 1470
rect 3640 1480 3690 1580
rect 3750 1860 3800 1970
rect 3750 1840 3760 1860
rect 3790 1840 3800 1860
rect 3750 1600 3800 1840
rect 3820 1860 3870 1910
rect 3820 1830 3830 1860
rect 3860 1830 3870 1860
rect 3820 1790 3870 1830
rect 3930 1860 3980 1880
rect 3930 1840 3940 1860
rect 3970 1840 3980 1860
rect 3750 1580 3760 1600
rect 3790 1580 3800 1600
rect 3750 1540 3800 1580
rect 3820 1600 3870 1660
rect 3820 1570 3830 1600
rect 3860 1570 3870 1600
rect 3820 1540 3870 1570
rect 3930 1600 3980 1840
rect 3930 1580 3940 1600
rect 3970 1580 3980 1600
rect 3930 1480 3980 1580
rect 4040 1870 4090 1960
rect 4040 1830 4050 1870
rect 4080 1830 4090 1870
rect 4040 1600 4090 1830
rect 4110 1860 4160 1910
rect 4110 1830 4120 1860
rect 4150 1830 4160 1860
rect 4110 1790 4160 1830
rect 5060 1860 5110 1880
rect 5060 1840 5070 1860
rect 5100 1840 5110 1860
rect 4040 1580 4050 1600
rect 4080 1580 4090 1600
rect 4040 1540 4090 1580
rect 4110 1600 4160 1660
rect 4110 1570 4120 1600
rect 4150 1570 4160 1600
rect 4110 1540 4160 1570
rect 5060 1600 5110 1840
rect 5060 1580 5070 1600
rect 5100 1580 5110 1600
rect 5060 1480 5110 1580
rect 5170 1860 5220 1970
rect 5170 1840 5180 1860
rect 5210 1840 5220 1860
rect 5170 1600 5220 1840
rect 5240 1860 5290 1910
rect 5240 1830 5250 1860
rect 5280 1830 5290 1860
rect 5240 1790 5290 1830
rect 5340 1860 5390 1880
rect 5340 1840 5350 1860
rect 5380 1840 5390 1860
rect 5170 1580 5180 1600
rect 5210 1580 5220 1600
rect 5170 1540 5220 1580
rect 5240 1600 5290 1660
rect 5240 1570 5250 1600
rect 5280 1570 5290 1600
rect 5240 1540 5290 1570
rect 5340 1600 5390 1840
rect 5340 1580 5350 1600
rect 5380 1580 5390 1600
rect 5340 1480 5390 1580
rect 5450 1860 5500 1970
rect 6090 1930 6420 1960
rect 5450 1840 5460 1860
rect 5490 1840 5500 1860
rect 5450 1600 5500 1840
rect 5520 1870 5570 1910
rect 5520 1840 5530 1870
rect 5560 1840 5570 1870
rect 5520 1790 5570 1840
rect 5770 1870 5810 1900
rect 5800 1840 5810 1870
rect 5770 1800 5810 1840
rect 6090 1860 6140 1930
rect 6090 1840 6100 1860
rect 6130 1840 6140 1860
rect 6090 1730 6140 1840
rect 5840 1720 6140 1730
rect 5840 1700 5850 1720
rect 5870 1700 6140 1720
rect 5840 1690 6140 1700
rect 5450 1580 5460 1600
rect 5490 1580 5500 1600
rect 5450 1540 5500 1580
rect 5520 1600 5570 1660
rect 5520 1570 5530 1600
rect 5560 1570 5570 1600
rect 5520 1540 5570 1570
rect 5630 1600 5690 1660
rect 5630 1560 5640 1600
rect 5680 1560 5690 1600
rect 5630 1540 5690 1560
rect 6090 1600 6140 1690
rect 6090 1580 6100 1600
rect 6130 1580 6140 1600
rect 5960 1540 6000 1550
rect 3640 1460 3980 1480
rect 4700 1470 5390 1480
rect 4700 1440 4730 1470
rect 4790 1440 4870 1470
rect 4930 1440 5390 1470
rect 4700 1430 5390 1440
rect 5960 1520 5970 1540
rect 5990 1520 6000 1540
rect 6090 1530 6140 1580
rect 6200 1860 6250 1910
rect 6200 1840 6210 1860
rect 6240 1840 6250 1860
rect 6200 1600 6250 1840
rect 6270 1870 6320 1910
rect 6270 1840 6280 1870
rect 6310 1840 6320 1870
rect 6270 1790 6320 1840
rect 6370 1860 6420 1930
rect 6370 1840 6380 1860
rect 6410 1840 6420 1860
rect 6200 1580 6210 1600
rect 6240 1580 6250 1600
rect 5960 1410 6000 1520
rect 6200 1450 6250 1580
rect 6270 1600 6320 1660
rect 6270 1570 6280 1600
rect 6310 1570 6320 1600
rect 6270 1540 6320 1570
rect 6370 1600 6420 1840
rect 6370 1580 6380 1600
rect 6410 1580 6420 1600
rect 6370 1530 6420 1580
rect 6480 1860 6530 1920
rect 6480 1840 6490 1860
rect 6520 1840 6530 1860
rect 6480 1730 6530 1840
rect 6550 1870 6600 1910
rect 6550 1840 6560 1870
rect 6590 1840 6600 1870
rect 6550 1790 6600 1840
rect 6660 1860 6710 1880
rect 6660 1840 6670 1860
rect 6700 1840 6710 1860
rect 6660 1730 6710 1840
rect 6480 1690 6710 1730
rect 6480 1600 6530 1690
rect 6480 1580 6490 1600
rect 6520 1580 6530 1600
rect 6480 1540 6530 1580
rect 6550 1600 6600 1660
rect 6550 1570 6560 1600
rect 6590 1570 6600 1600
rect 6550 1540 6600 1570
rect 6660 1600 6710 1690
rect 6660 1580 6670 1600
rect 6700 1580 6710 1600
rect 6660 1490 6710 1580
rect 6770 1860 6820 1960
rect 6770 1840 6780 1860
rect 6810 1840 6820 1860
rect 6770 1600 6820 1840
rect 6840 1860 6890 1910
rect 6840 1830 6850 1860
rect 6880 1830 6890 1860
rect 6840 1790 6890 1830
rect 6940 1860 6990 1880
rect 6940 1840 6950 1860
rect 6980 1840 6990 1860
rect 6770 1580 6780 1600
rect 6810 1580 6820 1600
rect 6770 1540 6820 1580
rect 6840 1600 6890 1660
rect 6840 1570 6850 1600
rect 6880 1570 6890 1600
rect 6840 1540 6890 1570
rect 6940 1600 6990 1840
rect 6940 1580 6950 1600
rect 6980 1580 6990 1600
rect 6940 1490 6990 1580
rect 7050 1870 7100 1960
rect 7050 1840 7060 1870
rect 7090 1840 7100 1870
rect 7050 1600 7100 1840
rect 7120 1860 7170 1910
rect 7120 1830 7130 1860
rect 7160 1830 7170 1860
rect 7120 1790 7170 1830
rect 7230 1810 7320 1820
rect 7230 1770 7240 1810
rect 7260 1791 7320 1810
rect 7260 1771 7300 1791
rect 7317 1771 7320 1791
rect 7260 1770 7320 1771
rect 7230 1760 7320 1770
rect 7380 1810 7420 1990
rect 8070 1900 8730 1920
rect 7700 1854 7705 1890
rect 7733 1854 7740 1890
rect 7700 1850 7710 1854
rect 7730 1850 7740 1854
rect 7700 1840 7740 1850
rect 8070 1880 8340 1900
rect 8360 1880 8700 1900
rect 8720 1880 8730 1900
rect 8070 1870 8730 1880
rect 8070 1810 8130 1870
rect 8850 1861 8890 1920
rect 7380 1770 7390 1810
rect 7410 1770 7420 1810
rect 7580 1800 8130 1810
rect 7580 1790 8080 1800
rect 7230 1680 7270 1760
rect 7380 1740 7420 1770
rect 7510 1780 7550 1790
rect 7510 1749 7520 1780
rect 7546 1749 7550 1780
rect 7580 1770 7590 1790
rect 7610 1770 8080 1790
rect 8110 1770 8130 1800
rect 7580 1760 8130 1770
rect 7510 1740 7550 1749
rect 7330 1730 7420 1740
rect 7330 1710 7340 1730
rect 7360 1710 7420 1730
rect 7330 1700 7420 1710
rect 7850 1720 7990 1730
rect 7230 1661 7320 1680
rect 7050 1580 7060 1600
rect 7090 1580 7100 1600
rect 7050 1540 7100 1580
rect 7120 1600 7170 1660
rect 7230 1630 7234 1661
rect 7266 1650 7320 1661
rect 7266 1630 7300 1650
rect 7317 1630 7320 1650
rect 7230 1620 7320 1630
rect 7380 1670 7420 1680
rect 7380 1630 7390 1670
rect 7410 1630 7420 1670
rect 7850 1670 7860 1720
rect 7890 1690 7950 1720
rect 7980 1690 7990 1720
rect 7890 1680 7990 1690
rect 7890 1670 7900 1680
rect 7850 1660 7900 1670
rect 7940 1650 7990 1680
rect 8060 1650 8130 1760
rect 8180 1720 8240 1840
rect 8850 1830 8856 1861
rect 8884 1830 8890 1861
rect 8850 1820 8890 1830
rect 9040 1869 9080 1920
rect 9040 1825 9044 1869
rect 9074 1825 9080 1869
rect 8380 1810 8630 1820
rect 8380 1780 8390 1810
rect 8430 1780 8630 1810
rect 8670 1780 8680 1820
rect 9040 1810 9080 1825
rect 10040 1880 10090 1900
rect 10040 1860 10050 1880
rect 10080 1860 10090 1880
rect 8380 1770 8680 1780
rect 8740 1740 8800 1750
rect 8540 1720 8600 1740
rect 8180 1700 8320 1720
rect 8180 1660 8190 1700
rect 8230 1670 8270 1700
rect 8310 1670 8320 1700
rect 8230 1660 8320 1670
rect 8540 1670 8550 1720
rect 8590 1670 8600 1720
rect 8740 1700 8750 1740
rect 8790 1700 8800 1740
rect 8740 1690 8800 1700
rect 7380 1620 8050 1630
rect 8180 1620 8240 1660
rect 7120 1570 7130 1600
rect 7160 1570 7170 1600
rect 7120 1540 7170 1570
rect 7380 1600 8020 1620
rect 8040 1600 8050 1620
rect 7380 1590 8050 1600
rect 6660 1470 6990 1490
rect 7380 1450 7420 1590
rect 6200 1430 7420 1450
rect 7950 1490 7990 1495
rect 7950 1459 7959 1490
rect 7986 1459 7990 1490
rect 2940 1390 6000 1410
rect 7950 1380 7990 1459
rect 8010 1492 8050 1496
rect 8010 1474 8020 1492
rect 8040 1474 8050 1492
rect 8010 1430 8050 1474
rect 8110 1490 8150 1496
rect 8540 1490 8600 1670
rect 10040 1620 10090 1860
rect 10040 1600 10050 1620
rect 10080 1600 10090 1620
rect 10040 1500 10090 1600
rect 10150 1880 10200 1990
rect 10150 1860 10160 1880
rect 10190 1860 10200 1880
rect 10150 1620 10200 1860
rect 10220 1890 10270 1930
rect 10220 1860 10230 1890
rect 10260 1860 10270 1890
rect 10220 1810 10270 1860
rect 10320 1880 10370 1900
rect 10320 1860 10330 1880
rect 10360 1860 10370 1880
rect 10150 1600 10160 1620
rect 10190 1600 10200 1620
rect 10150 1560 10200 1600
rect 10220 1620 10270 1680
rect 10220 1590 10230 1620
rect 10260 1590 10270 1620
rect 10220 1560 10270 1590
rect 10320 1620 10370 1860
rect 10320 1600 10330 1620
rect 10360 1600 10370 1620
rect 10320 1500 10370 1600
rect 10430 1880 10480 1980
rect 10430 1860 10440 1880
rect 10470 1860 10480 1880
rect 10430 1620 10480 1860
rect 10500 1890 10550 1930
rect 10500 1860 10510 1890
rect 10540 1860 10550 1890
rect 10500 1810 10550 1860
rect 11080 1880 11130 1900
rect 11080 1860 11090 1880
rect 11120 1860 11130 1880
rect 11080 1750 11130 1860
rect 10820 1740 11130 1750
rect 10820 1720 10830 1740
rect 10850 1720 11130 1740
rect 10820 1710 11130 1720
rect 10430 1600 10440 1620
rect 10470 1600 10480 1620
rect 10430 1560 10480 1600
rect 10500 1620 10550 1680
rect 10500 1590 10510 1620
rect 10540 1590 10550 1620
rect 10500 1560 10550 1590
rect 10630 1610 10690 1670
rect 10630 1570 10640 1610
rect 10680 1570 10690 1610
rect 10630 1550 10690 1570
rect 10750 1600 10790 1640
rect 10750 1559 10755 1600
rect 10785 1559 10790 1600
rect 11080 1620 11130 1710
rect 11080 1600 11090 1620
rect 11120 1600 11130 1620
rect 10750 1510 10790 1559
rect 10940 1560 10980 1580
rect 10940 1530 10950 1560
rect 10970 1530 10980 1560
rect 8110 1470 8120 1490
rect 8140 1470 8600 1490
rect 8110 1460 8600 1470
rect 9640 1490 10370 1500
rect 9640 1450 9670 1490
rect 9730 1450 9810 1490
rect 9870 1450 10370 1490
rect 9640 1440 10370 1450
rect 8010 1410 8020 1430
rect 8040 1410 8050 1430
rect 10940 1410 10980 1530
rect 11080 1490 11130 1600
rect 11190 1880 11240 1930
rect 11190 1860 11200 1880
rect 11230 1860 11240 1880
rect 11190 1620 11240 1860
rect 11260 1900 11310 1930
rect 11260 1860 11270 1900
rect 11300 1860 11310 1900
rect 11260 1810 11310 1860
rect 11360 1880 11410 1900
rect 11360 1860 11370 1880
rect 11400 1860 11410 1880
rect 11190 1590 11200 1620
rect 11230 1590 11240 1620
rect 11190 1560 11240 1590
rect 11260 1620 11310 1680
rect 11260 1590 11270 1620
rect 11300 1590 11310 1620
rect 11260 1560 11310 1590
rect 11360 1620 11410 1860
rect 11360 1600 11370 1620
rect 11400 1600 11410 1620
rect 11360 1490 11410 1600
rect 11470 1880 11520 1940
rect 11470 1860 11480 1880
rect 11510 1860 11520 1880
rect 11470 1750 11520 1860
rect 11540 1890 11590 1930
rect 11540 1860 11550 1890
rect 11580 1860 11590 1890
rect 11540 1810 11590 1860
rect 11640 1880 11690 1900
rect 11640 1860 11650 1880
rect 11680 1860 11690 1880
rect 11640 1750 11690 1860
rect 11470 1710 11690 1750
rect 11470 1620 11520 1710
rect 11470 1600 11480 1620
rect 11510 1600 11520 1620
rect 11470 1560 11520 1600
rect 11540 1620 11590 1680
rect 11540 1590 11550 1620
rect 11580 1590 11590 1620
rect 11540 1560 11590 1590
rect 11640 1620 11690 1710
rect 11640 1600 11650 1620
rect 11680 1600 11690 1620
rect 11080 1440 11410 1490
rect 11640 1500 11690 1600
rect 11750 1880 11800 1980
rect 11750 1860 11760 1880
rect 11790 1860 11800 1880
rect 11750 1620 11800 1860
rect 11820 1880 11870 1930
rect 12040 1900 12090 1990
rect 11820 1850 11830 1880
rect 11860 1850 11870 1880
rect 11820 1810 11870 1850
rect 11930 1880 11980 1900
rect 11930 1860 11940 1880
rect 11970 1860 11980 1880
rect 11750 1600 11760 1620
rect 11790 1600 11800 1620
rect 11750 1560 11800 1600
rect 11820 1620 11870 1680
rect 11820 1590 11830 1620
rect 11860 1590 11870 1620
rect 11820 1560 11870 1590
rect 11930 1620 11980 1860
rect 11930 1600 11940 1620
rect 11970 1600 11980 1620
rect 11930 1500 11980 1600
rect 12040 1860 12050 1900
rect 12080 1860 12090 1900
rect 12040 1620 12090 1860
rect 12110 1880 12160 1930
rect 12110 1850 12120 1880
rect 12150 1850 12160 1880
rect 12110 1810 12160 1850
rect 12040 1600 12050 1620
rect 12080 1600 12090 1620
rect 12040 1560 12090 1600
rect 12110 1620 12160 1680
rect 12110 1590 12120 1620
rect 12150 1590 12160 1620
rect 12110 1560 12160 1590
rect 11640 1440 11980 1500
rect 8010 1390 10980 1410
<< via1 >>
rect 2230 1860 2260 1880
rect 2230 1850 2260 1860
rect 2230 1600 2260 1610
rect 2230 1580 2260 1600
rect 2510 1850 2540 1870
rect 2510 1840 2540 1850
rect 2754 1900 2787 1901
rect 2754 1880 2760 1900
rect 2760 1880 2780 1900
rect 2780 1880 2787 1900
rect 2754 1873 2787 1880
rect 2510 1590 2540 1600
rect 2510 1570 2540 1590
rect 2610 1570 2650 1600
rect 2610 1560 2650 1570
rect 3260 1840 3290 1860
rect 3260 1830 3290 1840
rect 3260 1590 3290 1600
rect 3260 1570 3290 1590
rect 3550 1840 3580 1860
rect 3550 1830 3580 1840
rect 3550 1590 3580 1600
rect 3550 1570 3580 1590
rect 3830 1840 3860 1860
rect 3830 1830 3860 1840
rect 3830 1590 3860 1600
rect 3830 1570 3860 1590
rect 4050 1860 4080 1870
rect 4050 1840 4080 1860
rect 4050 1830 4080 1840
rect 4120 1840 4150 1860
rect 4120 1830 4150 1840
rect 4120 1590 4150 1600
rect 4120 1570 4150 1590
rect 5250 1840 5280 1860
rect 5250 1830 5280 1840
rect 5250 1590 5280 1600
rect 5250 1570 5280 1590
rect 5530 1850 5560 1870
rect 5530 1840 5560 1850
rect 5770 1860 5800 1870
rect 5770 1840 5780 1860
rect 5780 1840 5800 1860
rect 5530 1590 5560 1600
rect 5530 1570 5560 1590
rect 5640 1570 5680 1600
rect 5640 1560 5680 1570
rect 6280 1850 6310 1870
rect 6280 1840 6310 1850
rect 6280 1590 6310 1600
rect 6280 1570 6310 1590
rect 6560 1850 6590 1870
rect 6560 1840 6590 1850
rect 6560 1590 6590 1600
rect 6560 1570 6590 1590
rect 6850 1840 6880 1860
rect 6850 1830 6880 1840
rect 6850 1590 6880 1600
rect 6850 1570 6880 1590
rect 7060 1860 7090 1870
rect 7060 1840 7090 1860
rect 7130 1840 7160 1860
rect 7130 1830 7160 1840
rect 7705 1880 7733 1890
rect 7705 1854 7710 1880
rect 7710 1854 7730 1880
rect 7730 1854 7733 1880
rect 7520 1770 7546 1780
rect 7520 1750 7540 1770
rect 7540 1750 7546 1770
rect 7520 1749 7546 1750
rect 7234 1650 7266 1661
rect 7234 1630 7240 1650
rect 7240 1630 7260 1650
rect 7260 1630 7266 1650
rect 7860 1700 7890 1720
rect 7860 1680 7890 1700
rect 7860 1670 7890 1680
rect 8856 1860 8884 1861
rect 8856 1840 8860 1860
rect 8860 1840 8880 1860
rect 8880 1840 8884 1860
rect 8856 1830 8884 1840
rect 9044 1860 9074 1869
rect 9044 1830 9050 1860
rect 9050 1830 9070 1860
rect 9070 1830 9074 1860
rect 9044 1825 9074 1830
rect 8630 1810 8670 1820
rect 8630 1780 8670 1810
rect 8190 1680 8230 1700
rect 8190 1660 8230 1680
rect 8550 1690 8590 1720
rect 8550 1670 8590 1690
rect 8750 1710 8790 1740
rect 8750 1700 8790 1710
rect 7130 1590 7160 1600
rect 7130 1570 7160 1590
rect 7959 1470 7960 1490
rect 7960 1470 7980 1490
rect 7980 1470 7986 1490
rect 7959 1459 7986 1470
rect 10230 1870 10260 1890
rect 10230 1860 10260 1870
rect 10230 1610 10260 1620
rect 10230 1590 10260 1610
rect 10510 1870 10540 1890
rect 10510 1860 10540 1870
rect 10510 1610 10540 1620
rect 10510 1590 10540 1610
rect 10640 1580 10680 1610
rect 10640 1570 10680 1580
rect 10755 1580 10785 1600
rect 10755 1560 10760 1580
rect 10760 1560 10780 1580
rect 10780 1560 10785 1580
rect 10755 1559 10785 1560
rect 11270 1890 11300 1900
rect 11270 1870 11300 1890
rect 11270 1860 11300 1870
rect 11200 1600 11230 1620
rect 11200 1590 11230 1600
rect 11270 1610 11300 1620
rect 11270 1590 11300 1610
rect 11550 1870 11580 1890
rect 11550 1860 11580 1870
rect 11550 1610 11580 1620
rect 11550 1590 11580 1610
rect 11830 1860 11860 1880
rect 11830 1850 11860 1860
rect 11830 1610 11860 1620
rect 11830 1590 11860 1610
rect 12050 1880 12080 1900
rect 12050 1860 12080 1880
rect 12120 1860 12150 1880
rect 12120 1850 12150 1860
rect 12120 1610 12150 1620
rect 12120 1590 12150 1610
<< metal2 >>
rect 1160 2000 12230 2020
rect 2230 1880 2260 2000
rect 2230 1840 2260 1850
rect 2510 1870 2540 2000
rect 2750 1901 2790 2000
rect 2750 1873 2754 1901
rect 2787 1873 2790 1901
rect 2750 1860 2790 1873
rect 3260 1860 3290 2000
rect 2510 1830 2540 1840
rect 3260 1820 3290 1830
rect 3550 1860 3580 2000
rect 3550 1820 3580 1830
rect 3830 1860 3860 2000
rect 3830 1820 3860 1830
rect 4050 1870 4080 2000
rect 4050 1820 4080 1830
rect 4120 1860 4150 2000
rect 4120 1820 4150 1830
rect 5250 1860 5280 2000
rect 5530 1880 5560 2000
rect 5530 1870 5810 1880
rect 5560 1840 5770 1870
rect 5800 1840 5810 1870
rect 5530 1830 5810 1840
rect 6280 1870 6310 2000
rect 6280 1830 6310 1840
rect 6560 1870 6590 2000
rect 6560 1830 6590 1840
rect 6850 1860 6880 2000
rect 7050 1870 7100 2000
rect 7050 1840 7060 1870
rect 7090 1840 7100 1870
rect 7050 1830 7100 1840
rect 7130 1860 7160 2000
rect 5250 1820 5280 1830
rect 6850 1820 6880 1830
rect 7130 1820 7160 1830
rect 7510 1780 7550 2000
rect 7700 1890 7740 2000
rect 7700 1854 7705 1890
rect 7733 1854 7740 1890
rect 7700 1840 7740 1854
rect 7510 1749 7520 1780
rect 7546 1749 7550 1780
rect 7510 1740 7550 1749
rect 7850 1720 7900 1730
rect 7850 1670 7860 1720
rect 7890 1670 7900 1720
rect 7230 1661 7270 1670
rect 2230 1610 2260 1620
rect 2230 1390 2260 1580
rect 2510 1600 2540 1610
rect 2510 1390 2540 1570
rect 2600 1600 2660 1660
rect 2600 1560 2610 1600
rect 2650 1560 2660 1600
rect 2600 1540 2660 1560
rect 3260 1600 3290 1610
rect 3260 1390 3290 1570
rect 3550 1600 3580 1610
rect 3550 1390 3580 1570
rect 3830 1600 3860 1610
rect 3830 1390 3860 1570
rect 4120 1600 4150 1610
rect 4120 1390 4150 1570
rect 5250 1600 5280 1610
rect 5250 1390 5280 1570
rect 5530 1600 5560 1610
rect 5530 1390 5560 1570
rect 5630 1600 5690 1660
rect 7230 1630 7234 1661
rect 7266 1630 7270 1661
rect 5630 1560 5640 1600
rect 5680 1560 5690 1600
rect 5630 1540 5690 1560
rect 6280 1600 6310 1610
rect 6280 1390 6310 1570
rect 6560 1600 6590 1610
rect 6560 1390 6590 1570
rect 6850 1600 6880 1610
rect 6850 1390 6880 1570
rect 7130 1600 7160 1610
rect 7130 1390 7160 1570
rect 7230 1390 7270 1630
rect 7850 1390 7900 1670
rect 8180 1700 8240 1730
rect 8180 1660 8190 1700
rect 8230 1660 8240 1700
rect 8550 1720 8590 2000
rect 8620 1820 8680 1970
rect 8620 1780 8630 1820
rect 8670 1780 8680 1820
rect 8620 1770 8680 1780
rect 8740 1740 8800 2000
rect 8850 1861 8890 2000
rect 8850 1830 8856 1861
rect 8884 1830 8890 1861
rect 8850 1810 8890 1830
rect 9040 1869 9080 2000
rect 9040 1825 9044 1869
rect 9074 1825 9080 1869
rect 10230 1890 10260 2000
rect 10230 1850 10260 1860
rect 10510 1890 10540 2000
rect 10510 1850 10540 1860
rect 11270 1900 11300 2000
rect 11270 1850 11300 1860
rect 11550 1890 11580 2000
rect 11550 1850 11580 1860
rect 11830 1880 11860 2000
rect 11830 1830 11860 1850
rect 12040 1900 12090 2000
rect 12040 1860 12050 1900
rect 12080 1860 12090 1900
rect 9040 1810 9080 1825
rect 12040 1820 12090 1860
rect 12120 1880 12150 2000
rect 12120 1820 12150 1850
rect 8740 1700 8750 1740
rect 8790 1700 8800 1740
rect 8740 1690 8800 1700
rect 8550 1660 8590 1670
rect 7950 1490 7990 1495
rect 7950 1459 7959 1490
rect 7986 1459 7990 1490
rect 7950 1390 7990 1459
rect 8180 1390 8240 1660
rect 10230 1620 10260 1630
rect 10230 1390 10260 1590
rect 10510 1620 10540 1630
rect 10510 1390 10540 1590
rect 10630 1610 10690 1670
rect 10630 1570 10640 1610
rect 10680 1570 10690 1610
rect 10630 1550 10690 1570
rect 10750 1600 10790 1640
rect 10750 1559 10755 1600
rect 10785 1559 10790 1600
rect 10750 1390 10790 1559
rect 11190 1620 11240 1640
rect 11190 1590 11200 1620
rect 11230 1590 11240 1620
rect 11190 1390 11240 1590
rect 11270 1620 11300 1630
rect 11270 1390 11300 1590
rect 11550 1620 11580 1630
rect 11550 1390 11580 1590
rect 11830 1620 11860 1630
rect 11830 1390 11860 1590
rect 12120 1620 12150 1630
rect 12120 1390 12150 1590
rect 1150 1370 12190 1390
<< labels >>
flabel metal2 1280 2000 1310 2010 1 FreeSans 80 0 0 0 VDD
port 1 n
flabel metal2 1340 1370 1370 1380 1 FreeSans 80 0 0 0 GND
port 2 n
flabel metal1 2150 1950 2200 1970 1 FreeSans 80 0 0 0 VX
port 6 n
flabel metal1 2440 1950 2470 1960 1 FreeSans 80 0 0 0 CA0
port 4 n
flabel pmos 2880 1740 2920 1760 1 FreeSans 80 0 0 0 M4
flabel metal1 3760 1950 3790 1960 1 FreeSans 80 0 0 0 Vd
port 8 n
flabel metal1 3180 1700 3230 1720 1 FreeSans 80 0 0 0 M6Drain
flabel metal1 5180 1950 5210 1960 1 FreeSans 80 0 0 0 VFS2
port 9 n
flabel metal1 5460 1950 5490 1960 1 FreeSans 80 0 0 0 CA1
port 10 n
flabel pmos 5900 1740 5940 1760 1 FreeSans 80 0 0 0 M5
flabel metal1 6210 1700 6240 1710 1 FreeSans 80 0 0 0 M7Drain
flabel metal1 6780 1940 6810 1950 1 FreeSans 80 0 0 0 Vd
flabel nmos 7330 1780 7370 1810 1 FreeSans 80 0 0 0 M6
flabel nmos 7330 1640 7370 1670 1 FreeSans 80 0 0 0 M7
flabel pmos 7640 1730 7680 1750 1 FreeSans 80 0 0 0 M9
flabel pmos 8060 1470 8100 1490 1 FreeSans 80 0 0 0 M2
flabel nmos 8010 1730 8050 1750 1 FreeSans 80 0 0 0 M8
flabel nmos 8330 1740 8370 1760 1 FreeSans 80 0 0 0 M11
flabel pmos 8690 1730 8730 1750 1 FreeSans 80 0 0 0 M10
flabel pmos 8980 1710 9020 1730 1 FreeSans 80 0 0 0 M3
flabel metal2 8630 1930 8670 1940 1 FreeSans 80 0 0 0 bj
port 11 n
flabel metal1 10150 1960 10200 1980 1 FreeSans 80 0 0 0 Vbias
port 12 n
flabel metal1 10440 1960 10470 1970 1 FreeSans 80 0 0 0 CA2
port 13 n
flabel nmos 10880 1770 10920 1790 1 FreeSans 80 0 0 0 M1
flabel metal2 10630 1630 10690 1650 1 FreeSans 80 0 0 0 Vtun2
port 14 n
flabel metal2 5630 1620 5690 1640 1 FreeSans 80 0 0 0 Vtun1
port 15 n
flabel metal2 2600 1620 2660 1640 1 FreeSans 80 0 0 0 Vtun0
port 16 n
flabel metal1 11760 1960 11790 1970 1 FreeSans 80 0 0 0 Vd
port 8 n
<< end >>
