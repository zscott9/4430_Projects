* SPICE3 file created from sky130_hilas_Bootstrap01.ext - technology: sky130A

.option scale=10000u

.subckt sky130_hilas_Bootstrap01 RESIST VPWR VGND PBIAS NBIAS
X0 NBIAS PBIAS VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=581 l=20
X1 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X2 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X3 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X4 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X5 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X6 VPWR PBIAS PBIAS VPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=581 l=20
X7 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X8 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X9 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X10 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
R0 a_n535_n59# a_n454_n612# sky130_fd_pr__res_generic_po w=42 l=507
X11 NBIAS NBIAS VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=200 l=20
R1 RESIST a_n535_n59# sky130_fd_pr__res_generic_po w=42 l=507
X12 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X13 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X14 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X15 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X16 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X17 PBIAS NBIAS a_n454_n612# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
X18 a_n454_n612# NBIAS PBIAS VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=596 l=20
C0 PBIAS a_n454_n612# 15.95fF
.ends
