magic
tech sky130A
timestamp 1699313461
<< nwell >>
rect 0 300 3690 610
<< psubdiff >>
rect 0 110 70 130
rect 0 70 10 110
rect 50 70 70 110
rect 0 50 70 70
<< nsubdiff >>
rect 30 580 110 590
rect 30 540 50 580
rect 90 540 110 580
rect 30 520 110 540
<< psubdiffcont >>
rect 10 70 50 110
<< nsubdiffcont >>
rect 50 540 90 580
<< locali >>
rect 50 590 90 600
rect 40 580 60 590
rect 80 580 100 590
rect 40 540 50 580
rect 90 540 100 580
rect 40 530 100 540
rect 0 110 60 120
rect 0 70 10 110
rect 50 70 60 110
rect 0 60 60 70
<< viali >>
rect 60 580 80 590
rect 60 570 80 580
rect 20 70 40 90
<< metal1 >>
rect 50 600 100 610
rect 50 570 60 600
rect 90 570 100 600
rect 50 560 100 570
rect 10 100 60 110
rect 10 70 20 100
rect 50 70 60 100
rect 10 60 60 70
<< via1 >>
rect 60 590 90 600
rect 60 570 80 590
rect 80 570 90 590
rect 20 90 50 100
rect 20 70 40 90
rect 40 70 50 90
<< metal2 >>
rect 0 610 3690 650
rect 50 600 100 610
rect 50 570 60 600
rect 90 570 100 600
rect 50 560 100 570
rect 10 100 60 110
rect 10 70 20 100
rect 50 70 60 100
rect 10 40 60 70
rect 0 0 3690 40
<< labels >>
rlabel metal2 0 610 20 650 1 vdd
port 1 n
<< end >>
