magic
tech sky130A
timestamp 1697497807
<< nwell >>
rect 0 210 520 590
rect 0 50 1400 210
<< nmos >>
rect 610 450 650 530
rect 790 439 830 530
rect 970 440 1010 580
rect 1060 480 1100 530
rect 610 280 650 360
rect 790 280 830 360
rect 880 280 920 360
rect 1060 280 1100 360
rect 1150 290 1190 340
<< pmos >>
rect 90 80 130 240
rect 270 80 310 560
rect 360 80 400 560
rect 540 80 580 160
rect 630 80 670 160
rect 720 82 760 160
rect 950 90 990 140
rect 1040 90 1080 140
rect 1210 70 1250 150
rect 1300 70 1340 150
<< ndiff >>
rect 920 570 970 580
rect 560 520 610 530
rect 560 460 570 520
rect 600 460 610 520
rect 560 450 610 460
rect 650 520 700 530
rect 650 460 660 520
rect 690 460 700 520
rect 650 450 700 460
rect 740 520 790 530
rect 740 450 750 520
rect 780 450 790 520
rect 740 439 790 450
rect 830 520 880 530
rect 830 450 840 520
rect 870 450 880 520
rect 830 439 880 450
rect 920 450 930 570
rect 960 450 970 570
rect 920 440 970 450
rect 1010 530 1040 580
rect 1010 520 1060 530
rect 1010 490 1020 520
rect 1050 490 1060 520
rect 1010 480 1060 490
rect 1100 520 1150 530
rect 1100 490 1110 520
rect 1140 490 1150 520
rect 1100 480 1150 490
rect 1010 440 1040 480
rect 560 350 610 360
rect 560 290 570 350
rect 600 290 610 350
rect 560 280 610 290
rect 650 350 700 360
rect 650 290 660 350
rect 690 290 700 350
rect 650 280 700 290
rect 740 350 790 360
rect 740 290 750 350
rect 780 290 790 350
rect 740 280 790 290
rect 830 350 880 360
rect 830 290 840 350
rect 870 290 880 350
rect 830 280 880 290
rect 920 350 970 360
rect 920 290 930 350
rect 960 290 970 350
rect 920 280 970 290
rect 1010 350 1060 360
rect 1010 290 1020 350
rect 1050 290 1060 350
rect 1010 280 1060 290
rect 1100 340 1140 360
rect 1100 330 1150 340
rect 1100 300 1110 330
rect 1140 300 1150 330
rect 1100 290 1150 300
rect 1190 330 1240 340
rect 1190 300 1200 330
rect 1230 300 1240 330
rect 1190 290 1240 300
rect 1100 280 1140 290
<< pdiff >>
rect 220 550 270 560
rect 40 230 90 240
rect 40 90 50 230
rect 80 90 90 230
rect 40 80 90 90
rect 130 230 180 240
rect 130 90 140 230
rect 170 90 180 230
rect 130 80 180 90
rect 220 90 230 550
rect 260 90 270 550
rect 220 80 270 90
rect 310 550 360 560
rect 310 90 320 550
rect 350 90 360 550
rect 310 80 360 90
rect 400 550 450 560
rect 400 90 410 550
rect 440 90 450 550
rect 400 80 450 90
rect 490 150 540 160
rect 490 90 500 150
rect 530 90 540 150
rect 490 80 540 90
rect 580 130 630 160
rect 580 100 590 130
rect 620 100 630 130
rect 580 80 630 100
rect 670 82 720 160
rect 760 140 810 160
rect 1160 140 1210 150
rect 760 100 770 140
rect 800 100 810 140
rect 760 82 810 100
rect 900 130 950 140
rect 900 100 910 130
rect 940 100 950 130
rect 900 90 950 100
rect 990 130 1040 140
rect 990 100 1000 130
rect 1030 100 1040 130
rect 990 90 1040 100
rect 1080 130 1130 140
rect 1080 100 1090 130
rect 1120 100 1130 130
rect 1080 90 1130 100
rect 670 80 700 82
rect 790 80 810 82
rect 1160 80 1170 140
rect 1200 80 1210 140
rect 1160 70 1210 80
rect 1250 130 1300 150
rect 1250 90 1260 130
rect 1290 90 1300 130
rect 1250 70 1300 90
rect 1340 140 1380 150
rect 1340 80 1350 140
rect 1370 80 1380 140
rect 1340 70 1380 80
<< ndiffc >>
rect 570 460 600 520
rect 660 460 690 520
rect 750 450 780 520
rect 840 450 870 520
rect 930 450 960 570
rect 1020 490 1050 520
rect 1110 490 1140 520
rect 570 290 600 350
rect 660 290 690 350
rect 750 290 780 350
rect 840 290 870 350
rect 930 290 960 350
rect 1020 290 1050 350
rect 1110 300 1140 330
rect 1200 300 1230 330
<< pdiffc >>
rect 50 90 80 230
rect 140 90 170 230
rect 230 90 260 550
rect 320 90 350 550
rect 410 90 440 550
rect 500 90 530 150
rect 590 100 620 130
rect 770 100 800 140
rect 910 100 940 130
rect 1000 100 1030 130
rect 1090 100 1120 130
rect 1170 80 1200 140
rect 1260 90 1290 130
rect 1350 80 1370 140
<< psubdiff >>
rect 1310 490 1390 500
rect 1310 390 1330 490
rect 1370 390 1390 490
rect 1310 370 1390 390
<< nsubdiff >>
rect 40 530 170 570
rect 40 400 80 530
rect 130 400 170 530
rect 40 360 170 400
<< psubdiffcont >>
rect 1330 390 1370 490
<< nsubdiffcont >>
rect 80 400 130 530
<< poly >>
rect 270 610 310 620
rect 270 590 280 610
rect 300 590 310 610
rect 270 560 310 590
rect 360 610 400 620
rect 360 590 370 610
rect 390 590 400 610
rect 360 560 400 590
rect 610 580 650 590
rect 970 580 1010 600
rect 1060 590 1100 600
rect 610 560 620 580
rect 640 560 650 580
rect 90 290 130 300
rect 90 270 100 290
rect 120 270 130 290
rect 90 240 130 270
rect 610 530 650 560
rect 740 570 830 580
rect 740 550 750 570
rect 800 550 830 570
rect 740 540 830 550
rect 790 530 830 540
rect 610 360 650 450
rect 1060 560 1070 590
rect 1090 560 1100 590
rect 1060 530 1100 560
rect 790 420 830 439
rect 970 410 1010 440
rect 970 390 980 410
rect 1000 390 1010 410
rect 970 380 1010 390
rect 790 360 830 380
rect 880 360 920 380
rect 1060 360 1100 480
rect 1150 340 1190 360
rect 610 250 650 280
rect 790 250 830 280
rect 790 230 800 250
rect 820 230 830 250
rect 790 220 830 230
rect 880 250 920 280
rect 1060 260 1100 280
rect 1150 270 1190 290
rect 1150 260 1240 270
rect 880 230 890 250
rect 910 230 920 250
rect 1150 240 1200 260
rect 1230 240 1240 260
rect 1150 230 1240 240
rect 1300 230 1380 240
rect 880 220 920 230
rect 540 210 580 220
rect 540 190 550 210
rect 570 190 580 210
rect 1300 210 1330 230
rect 1370 210 1380 230
rect 1300 200 1380 210
rect 540 160 580 190
rect 630 160 670 180
rect 720 160 760 180
rect 950 140 990 160
rect 1040 140 1080 160
rect 1210 150 1250 200
rect 1300 150 1340 200
rect 90 60 130 80
rect 270 60 310 80
rect 360 60 400 80
rect 540 60 580 80
rect 630 60 670 80
rect 540 40 670 60
rect 720 50 760 82
rect 720 20 730 50
rect 750 20 760 50
rect 950 70 990 90
rect 950 60 1000 70
rect 950 40 970 60
rect 990 40 1000 60
rect 950 30 1000 40
rect 1040 60 1080 90
rect 1210 60 1250 70
rect 1040 50 1250 60
rect 1300 50 1340 70
rect 1040 30 1100 50
rect 1130 30 1250 50
rect 1040 20 1250 30
rect 720 10 760 20
<< polycont >>
rect 280 590 300 610
rect 370 590 390 610
rect 620 560 640 580
rect 100 270 120 290
rect 750 550 800 570
rect 1070 560 1090 590
rect 980 390 1000 410
rect 800 230 820 250
rect 890 230 910 250
rect 1200 240 1230 260
rect 550 190 570 210
rect 1330 210 1370 230
rect 730 20 750 50
rect 970 40 990 60
rect 1100 30 1130 50
<< locali >>
rect 270 610 310 620
rect 270 590 280 610
rect 300 590 310 610
rect 270 580 310 590
rect 360 610 400 620
rect 360 590 370 610
rect 390 590 400 610
rect 1060 590 1100 600
rect 360 580 400 590
rect 610 580 700 590
rect 610 560 620 580
rect 640 560 700 580
rect 220 550 270 560
rect 70 530 90 550
rect 120 530 140 550
rect 70 400 80 530
rect 130 400 140 530
rect 70 390 140 400
rect 90 290 130 300
rect 90 270 100 290
rect 120 270 130 290
rect 90 260 130 270
rect 40 230 90 240
rect 40 90 50 230
rect 80 90 90 230
rect 40 80 90 90
rect 130 230 180 240
rect 130 90 140 230
rect 170 90 180 230
rect 130 80 180 90
rect 220 90 230 550
rect 260 90 270 550
rect 220 80 270 90
rect 310 550 360 560
rect 310 90 320 550
rect 350 90 360 550
rect 310 80 360 90
rect 400 550 450 560
rect 610 550 700 560
rect 400 90 410 550
rect 440 90 450 550
rect 660 530 700 550
rect 740 570 810 580
rect 740 550 750 570
rect 800 550 810 570
rect 740 540 760 550
rect 790 540 810 550
rect 920 570 970 580
rect 560 520 610 530
rect 560 460 570 520
rect 600 460 610 520
rect 560 350 610 460
rect 650 520 700 530
rect 830 520 880 530
rect 650 460 660 520
rect 690 460 700 520
rect 650 450 700 460
rect 740 450 750 520
rect 780 450 790 520
rect 740 439 790 450
rect 830 450 840 520
rect 870 450 880 520
rect 830 440 880 450
rect 920 450 930 570
rect 960 450 970 570
rect 1060 560 1070 590
rect 1090 560 1100 590
rect 1060 550 1100 560
rect 1010 520 1060 530
rect 1010 490 1020 520
rect 1050 490 1060 520
rect 1010 480 1060 490
rect 1100 520 1150 530
rect 1100 490 1110 520
rect 1140 490 1150 520
rect 1100 480 1150 490
rect 1310 490 1390 510
rect 920 440 970 450
rect 970 410 1010 420
rect 970 390 980 410
rect 1000 390 1010 410
rect 970 380 1010 390
rect 1310 390 1330 490
rect 1370 390 1390 490
rect 1310 370 1390 390
rect 560 290 570 350
rect 600 290 610 350
rect 560 280 610 290
rect 650 350 700 360
rect 650 290 660 350
rect 690 290 700 350
rect 650 280 700 290
rect 740 350 790 360
rect 740 290 750 350
rect 780 290 790 350
rect 740 260 790 290
rect 830 350 880 360
rect 830 290 840 350
rect 870 290 880 350
rect 830 280 880 290
rect 920 350 970 360
rect 920 290 930 350
rect 960 290 970 350
rect 920 280 970 290
rect 1010 350 1060 360
rect 1010 290 1020 350
rect 1050 290 1060 350
rect 1100 330 1150 340
rect 1100 300 1110 330
rect 1140 300 1150 330
rect 1100 290 1150 300
rect 1190 330 1240 340
rect 1190 300 1200 330
rect 1230 300 1240 330
rect 1190 290 1240 300
rect 1010 280 1060 290
rect 740 230 750 260
rect 780 250 920 260
rect 780 230 800 250
rect 820 230 890 250
rect 910 230 920 250
rect 740 220 920 230
rect 540 210 580 220
rect 540 200 550 210
rect 400 80 450 90
rect 490 190 550 200
rect 570 200 580 210
rect 940 200 970 280
rect 1020 260 1050 280
rect 1190 260 1240 270
rect 1020 230 1110 260
rect 1140 230 1150 260
rect 1190 240 1200 260
rect 1230 240 1240 260
rect 1190 230 1240 240
rect 1200 200 1240 230
rect 1320 240 1380 250
rect 1320 230 1340 240
rect 1320 210 1330 230
rect 1370 210 1380 240
rect 1320 200 1380 210
rect 570 190 970 200
rect 490 170 970 190
rect 1000 180 1010 200
rect 490 150 540 170
rect 490 90 500 150
rect 530 90 540 150
rect 760 140 810 150
rect 1000 140 1030 180
rect 1200 170 1300 200
rect 1160 140 1210 150
rect 590 130 620 140
rect 590 90 620 100
rect 760 100 770 140
rect 800 100 810 140
rect 760 90 810 100
rect 900 130 950 140
rect 900 100 910 130
rect 940 100 950 130
rect 900 90 950 100
rect 990 130 1040 140
rect 990 100 1000 130
rect 1030 100 1040 130
rect 990 90 1040 100
rect 1080 130 1130 140
rect 1080 100 1090 130
rect 1120 100 1130 130
rect 1080 90 1130 100
rect 490 80 540 90
rect 1160 80 1170 140
rect 1200 80 1210 140
rect 1250 130 1300 170
rect 1250 90 1260 130
rect 1290 90 1300 130
rect 1250 80 1300 90
rect 1340 140 1380 150
rect 1340 80 1350 140
rect 1370 80 1380 140
rect 950 60 1000 70
rect 400 50 760 60
rect 400 20 410 50
rect 440 20 730 50
rect 750 20 760 50
rect 950 40 970 60
rect 990 40 1000 60
rect 1030 50 1040 70
rect 1410 60 1450 70
rect 1090 50 1450 60
rect 950 30 1000 40
rect 1090 30 1100 50
rect 1130 30 1420 50
rect 1440 30 1450 50
rect 1090 20 1450 30
rect 400 10 760 20
<< viali >>
rect 280 590 300 610
rect 370 590 390 610
rect 620 560 640 580
rect 90 530 120 550
rect 100 270 120 290
rect 50 140 80 170
rect 140 90 170 120
rect 230 480 260 510
rect 320 90 350 120
rect 410 180 440 210
rect 760 550 790 570
rect 760 540 790 550
rect 660 470 690 500
rect 750 450 780 480
rect 840 450 870 520
rect 930 540 960 570
rect 1070 560 1090 590
rect 1020 490 1050 520
rect 1110 490 1140 520
rect 980 390 1000 410
rect 1340 430 1360 460
rect 570 320 600 350
rect 660 300 690 330
rect 840 290 870 320
rect 1110 300 1140 330
rect 1200 300 1230 330
rect 750 230 780 260
rect 1110 230 1140 260
rect 1340 230 1370 240
rect 1340 210 1370 230
rect 1010 180 1030 200
rect 500 90 530 120
rect 590 100 620 130
rect 770 100 800 140
rect 910 100 940 130
rect 1090 100 1120 130
rect 1170 90 1200 120
rect 1350 80 1370 110
rect 410 20 440 50
rect 1000 50 1030 70
rect 1420 30 1440 50
<< metal1 >>
rect 920 640 970 650
rect 80 610 90 640
rect 120 610 130 640
rect 270 610 310 620
rect 360 610 400 620
rect 80 550 130 610
rect 240 590 280 610
rect 300 590 310 610
rect 330 590 370 610
rect 390 590 400 610
rect 920 610 930 640
rect 960 610 970 640
rect 270 580 310 590
rect 360 580 400 590
rect 610 580 650 590
rect 610 560 620 580
rect 640 560 650 580
rect 610 550 650 560
rect 750 570 800 580
rect 80 530 90 550
rect 120 530 130 550
rect 750 540 760 570
rect 790 540 800 570
rect 750 530 800 540
rect 920 570 970 610
rect 920 540 930 570
rect 960 540 970 570
rect 1060 590 1100 600
rect 1060 560 1070 590
rect 1090 560 1100 590
rect 1060 550 1100 560
rect 920 530 970 540
rect 80 520 130 530
rect 660 520 710 530
rect 220 510 710 520
rect 220 480 230 510
rect 260 500 710 510
rect 260 480 660 500
rect 220 470 660 480
rect 690 470 710 500
rect 830 520 880 530
rect 650 460 710 470
rect 740 480 790 490
rect 740 450 750 480
rect 780 450 790 480
rect 740 420 790 450
rect 830 450 840 520
rect 870 450 880 520
rect 1010 520 1060 530
rect 1010 490 1020 520
rect 1050 490 1060 520
rect 1010 480 1060 490
rect 1100 520 1150 530
rect 1100 490 1110 520
rect 1140 490 1370 520
rect 1100 480 1150 490
rect 830 440 880 450
rect 1330 460 1370 490
rect 1100 430 1220 440
rect 650 380 790 420
rect 970 410 1040 420
rect 970 390 980 410
rect 1000 390 1040 410
rect 970 380 1040 390
rect 560 350 610 360
rect 560 320 570 350
rect 600 320 610 350
rect 500 310 540 320
rect 560 310 610 320
rect 650 330 710 380
rect 110 300 200 310
rect 50 290 160 300
rect 50 270 100 290
rect 120 270 160 290
rect 190 270 200 300
rect 50 260 200 270
rect 530 280 540 310
rect 650 300 660 330
rect 690 300 710 330
rect 740 330 750 360
rect 780 340 790 360
rect 780 330 880 340
rect 740 320 880 330
rect 740 310 790 320
rect 650 280 710 300
rect 830 290 840 320
rect 870 290 880 320
rect 500 250 540 280
rect 740 260 790 270
rect 400 210 450 220
rect 500 210 630 250
rect 400 180 410 210
rect 440 180 450 210
rect 40 170 90 180
rect 400 170 450 180
rect 40 140 50 170
rect 80 140 90 170
rect 40 130 90 140
rect 580 130 630 210
rect 740 230 750 260
rect 780 230 790 260
rect 740 210 790 230
rect 740 180 750 210
rect 780 180 790 210
rect 740 170 790 180
rect 130 120 360 130
rect 130 90 140 120
rect 170 90 320 120
rect 350 90 360 120
rect 490 120 540 130
rect 130 80 360 90
rect 400 100 450 110
rect 400 70 410 100
rect 440 70 450 100
rect 490 90 500 120
rect 530 90 540 120
rect 580 100 590 130
rect 620 100 630 130
rect 580 90 630 100
rect 760 140 810 150
rect 760 100 770 140
rect 800 100 810 140
rect 760 90 810 100
rect 490 80 540 90
rect 400 50 450 70
rect 400 20 410 50
rect 440 20 450 50
rect 400 10 450 20
rect 830 40 880 290
rect 1000 200 1040 380
rect 1100 400 1180 430
rect 1210 400 1220 430
rect 1330 430 1340 460
rect 1360 430 1370 460
rect 1330 420 1370 430
rect 1100 390 1220 400
rect 1100 330 1150 390
rect 1100 300 1110 330
rect 1140 300 1150 330
rect 1100 290 1150 300
rect 1190 330 1240 340
rect 1190 300 1200 330
rect 1230 300 1240 330
rect 1190 290 1240 300
rect 1100 260 1150 270
rect 1100 230 1110 260
rect 1140 230 1150 260
rect 1100 220 1150 230
rect 1330 240 1380 250
rect 1330 210 1340 240
rect 1370 210 1380 240
rect 1330 200 1380 210
rect 1000 180 1010 200
rect 1030 180 1040 200
rect 1250 190 1300 200
rect 1000 170 1040 180
rect 1080 160 1260 190
rect 1290 160 1300 190
rect 990 140 1040 150
rect 830 10 840 40
rect 870 10 880 40
rect 830 0 880 10
rect 900 130 950 140
rect 900 100 910 130
rect 940 100 950 130
rect 900 40 950 100
rect 990 110 1000 140
rect 1030 110 1040 140
rect 990 70 1040 110
rect 1080 130 1130 160
rect 1250 150 1300 160
rect 1080 100 1090 130
rect 1120 100 1130 130
rect 1080 90 1130 100
rect 1160 120 1210 130
rect 1160 90 1170 120
rect 1200 90 1210 120
rect 1160 80 1210 90
rect 1340 110 1380 120
rect 1340 80 1350 110
rect 1370 80 1380 110
rect 990 50 1000 70
rect 1030 50 1040 70
rect 990 40 1040 50
rect 1340 40 1380 80
rect 900 10 910 40
rect 940 10 950 40
rect 900 0 950 10
rect 1340 10 1350 40
rect 1410 110 1460 120
rect 1410 80 1420 110
rect 1450 80 1460 110
rect 1410 50 1460 80
rect 1410 30 1420 50
rect 1440 30 1460 50
rect 1410 20 1460 30
rect 1340 0 1380 10
<< via1 >>
rect 90 610 120 640
rect 930 610 960 640
rect 760 540 790 570
rect 660 470 690 500
rect 840 450 870 520
rect 1020 490 1050 520
rect 1110 490 1140 520
rect 570 320 600 350
rect 160 270 190 300
rect 500 280 530 310
rect 750 330 780 360
rect 410 180 440 210
rect 50 140 80 170
rect 750 180 780 210
rect 410 70 440 100
rect 500 90 530 120
rect 770 100 800 140
rect 1180 400 1210 430
rect 1200 300 1230 330
rect 1110 230 1140 260
rect 1340 210 1370 240
rect 1260 160 1290 190
rect 840 10 870 40
rect 1000 110 1030 140
rect 1170 90 1200 120
rect 910 10 940 40
rect 1350 10 1380 40
rect 1420 80 1450 110
<< metal2 >>
rect 0 640 1400 650
rect 0 610 90 640
rect 120 610 930 640
rect 960 610 1400 640
rect 50 180 80 610
rect 500 310 530 610
rect 750 570 800 580
rect 750 540 760 570
rect 790 540 800 570
rect 650 500 710 540
rect 750 530 800 540
rect 650 470 660 500
rect 690 470 710 500
rect 650 460 710 470
rect 830 520 880 570
rect 830 450 840 520
rect 870 450 880 520
rect 1010 520 1080 530
rect 1010 490 1020 520
rect 1070 490 1080 520
rect 1010 480 1080 490
rect 1100 520 1150 530
rect 1100 490 1110 520
rect 1140 490 1150 520
rect 560 350 750 360
rect 560 320 570 350
rect 600 330 750 350
rect 780 330 800 360
rect 600 320 800 330
rect 560 310 800 320
rect 150 300 200 310
rect 150 270 160 300
rect 190 270 200 300
rect 500 270 530 280
rect 150 260 200 270
rect 400 210 790 220
rect 400 180 410 210
rect 440 180 750 210
rect 780 180 790 210
rect 40 170 90 180
rect 400 170 790 180
rect 40 140 50 170
rect 80 140 90 170
rect 830 150 880 450
rect 1100 260 1150 490
rect 1170 430 1220 440
rect 1170 400 1180 430
rect 1210 400 1220 430
rect 1170 390 1220 400
rect 1250 340 1300 610
rect 1190 330 1300 340
rect 1190 300 1200 330
rect 1230 300 1300 330
rect 1190 290 1300 300
rect 1100 230 1110 260
rect 1140 230 1150 260
rect 40 130 90 140
rect 760 140 880 150
rect 490 120 540 130
rect 400 110 450 120
rect 400 70 410 110
rect 440 70 450 110
rect 490 90 500 120
rect 530 90 540 120
rect 760 100 770 140
rect 800 100 880 140
rect 990 140 1040 150
rect 1100 140 1150 230
rect 990 110 1000 140
rect 1030 110 1040 140
rect 990 100 1040 110
rect 760 90 880 100
rect 1080 90 1150 140
rect 1250 190 1300 290
rect 1330 240 1380 250
rect 1330 210 1340 240
rect 1370 210 1380 240
rect 1330 200 1380 210
rect 1250 160 1260 190
rect 1290 160 1300 190
rect 1250 130 1300 160
rect 490 80 540 90
rect 400 60 450 70
rect 1100 40 1150 90
rect 1170 120 1300 130
rect 1200 90 1300 120
rect 1170 80 1300 90
rect 1410 110 1460 120
rect 1410 80 1420 110
rect 1450 80 1460 110
rect 1410 70 1460 80
rect 0 10 840 40
rect 870 10 910 40
rect 940 10 1350 40
rect 1380 10 1460 40
rect 0 0 1460 10
<< via2 >>
rect 760 540 790 570
rect 660 470 690 500
rect 1040 490 1050 520
rect 1050 490 1070 520
rect 160 270 190 300
rect 1180 400 1210 430
rect 410 100 440 110
rect 410 80 440 100
rect 500 90 530 120
rect 1000 110 1030 140
rect 1340 210 1370 240
rect 1420 80 1450 110
<< metal3 >>
rect 750 570 840 590
rect 750 540 760 570
rect 790 540 840 570
rect 650 520 710 540
rect 750 530 840 540
rect 790 520 1080 530
rect 650 500 720 520
rect 650 470 660 500
rect 690 470 720 500
rect 790 490 1040 520
rect 1070 490 1080 520
rect 790 480 1080 490
rect 650 460 720 470
rect 670 360 720 460
rect 1160 440 1230 450
rect 1160 390 1170 440
rect 1220 390 1230 440
rect 1160 380 1230 390
rect 670 310 1040 360
rect 150 300 200 310
rect 50 270 160 300
rect 190 270 200 300
rect 50 260 200 270
rect 50 40 90 260
rect 490 120 950 160
rect 400 110 460 120
rect 400 70 410 110
rect 450 70 460 110
rect 490 90 500 120
rect 530 90 540 120
rect 490 70 540 90
rect 580 60 660 70
rect 580 40 600 60
rect 50 20 600 40
rect 640 20 660 60
rect 50 10 660 20
rect 900 50 950 120
rect 990 140 1040 310
rect 1330 240 1380 250
rect 990 110 1000 140
rect 1030 110 1040 140
rect 990 100 1040 110
rect 1300 210 1340 240
rect 1370 210 1380 240
rect 1300 170 1380 210
rect 1300 50 1340 170
rect 1410 120 1470 130
rect 1410 80 1420 120
rect 1460 80 1470 120
rect 1410 70 1470 80
rect 900 10 1340 50
rect 50 0 650 10
<< via3 >>
rect 1170 430 1220 440
rect 1170 400 1180 430
rect 1180 400 1210 430
rect 1210 400 1220 430
rect 1170 390 1220 400
rect 410 80 440 110
rect 440 80 450 110
rect 410 70 450 80
rect 600 20 640 60
rect 1420 110 1460 120
rect 1420 80 1450 110
rect 1450 80 1460 110
<< metal4 >>
rect 1160 440 1230 450
rect 1150 390 1170 440
rect 1220 390 1230 440
rect 1150 380 1230 390
rect 1150 270 1220 380
rect 400 220 1210 270
rect 400 110 460 220
rect 400 70 410 110
rect 450 70 460 110
rect 400 60 460 70
rect 580 120 1470 130
rect 580 80 1420 120
rect 1460 80 1470 120
rect 580 70 1470 80
rect 580 60 660 70
rect 580 20 600 60
rect 640 20 660 60
rect 580 10 660 20
<< labels >>
rlabel metal2 0 610 20 650 1 VDD
port 2 n
rlabel metal1 240 590 260 610 1 VIN1
port 3 n
rlabel metal1 330 590 350 610 1 VIN2
port 4 n
rlabel metal2 520 170 600 220 1 V26
rlabel metal1 740 380 790 420 1 V45
rlabel locali 940 210 970 260 1 V78
rlabel pdiff 670 82 720 160 1 V910
rlabel metal2 830 550 880 570 1 VOUT
port 6 n
rlabel metal1 50 260 100 300 1 PBIAS
port 7 n
rlabel ndiff 1010 480 1060 530 1 VCNACT
rlabel metal1 520 470 560 520 1 V13
rlabel pdiff 990 90 1040 140 1 VCNTEMP
rlabel metal1 1060 580 1100 600 1 NBIAS
port 8 n
rlabel pdiff 1250 70 1300 150 1 VCPTEMP
rlabel metal4 1160 380 1230 450 1 VCPACT
rlabel pdiffc 140 90 170 230 1 VINT
rlabel metal2 0 0 20 40 1 VGND
port 5 n
<< end >>
