** sch_path: /home/bard/4430_Projects/project2/sky130_hilas_Bootstrap01.sch
**.subckt sky130_hilas_Bootstrap01 VPWR NBIAS PBIAS VGND RESIST RESIST VPWR
*.iopin VPWR
*.iopin NBIAS
*.iopin PBIAS
*.iopin VGND
*.iopin RESIST
*.iopin RESIST
*.iopin VPWR
XM4 NBIAS NBIAS VGND VGND sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 NBIAS PBIAS VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.2 W=5.81 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 PBIAS NBIAS net1 VGND sky130_fd_pr__nfet_01v8 L=0.2 W=95.36 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 PBIAS PBIAS VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.2 W=5.81 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 RESIST net1 sky130_fd_pr__res_generic_po W=0.42 L=10.14 m=1
**.ends
.GLOBAL VGND
.end
