magic
tech sky130A
timestamp 1699375158
<< nwell >>
rect 0 40 1880 610
rect 3520 280 5200 610
rect 3520 40 4940 280
<< nmos >>
rect 2070 340 2370 540
rect 2870 340 3170 540
rect 5290 350 5590 550
rect 2070 100 2670 300
rect 2870 100 3470 300
rect 5010 140 5090 180
rect 5290 100 5590 300
<< pmos >>
rect 50 450 1850 550
rect 60 310 660 350
rect 3670 340 3970 540
rect 4160 340 4460 540
rect 4590 340 4890 540
rect 5060 360 5140 400
rect 40 110 1840 210
rect 3670 100 3970 300
rect 4160 100 4460 300
rect 4590 100 4890 300
<< ndiff >>
rect 2070 570 2370 580
rect 2070 550 2080 570
rect 2360 550 2370 570
rect 2070 540 2370 550
rect 2870 570 3170 580
rect 2870 550 2880 570
rect 3160 550 3170 570
rect 2870 540 3170 550
rect 5290 580 5590 590
rect 5290 560 5300 580
rect 5580 560 5590 580
rect 5290 550 5590 560
rect 2070 330 2370 340
rect 2870 330 3170 340
rect 2070 310 2080 330
rect 2360 310 2670 330
rect 2070 300 2670 310
rect 2870 310 2880 330
rect 3160 310 3470 330
rect 2870 300 3470 310
rect 5290 340 5590 350
rect 5290 310 5300 340
rect 5580 310 5590 340
rect 5290 300 5590 310
rect 5010 210 5090 220
rect 5010 190 5020 210
rect 5080 190 5090 210
rect 5010 180 5090 190
rect 5010 130 5090 140
rect 5010 110 5020 130
rect 5080 110 5090 130
rect 5010 100 5090 110
rect 2070 90 2670 100
rect 2070 70 2080 90
rect 2660 70 2670 90
rect 2070 60 2670 70
rect 2870 90 3470 100
rect 2870 70 2880 90
rect 3460 70 3470 90
rect 2870 60 3470 70
rect 5290 90 5590 100
rect 5290 70 5300 90
rect 5580 70 5590 90
rect 5290 60 5590 70
<< pdiff >>
rect 50 580 1850 590
rect 50 560 60 580
rect 1840 560 1850 580
rect 50 550 1850 560
rect 3670 570 3970 580
rect 3670 550 3680 570
rect 3960 550 3970 570
rect 3670 540 3970 550
rect 4160 570 4460 580
rect 4160 550 4170 570
rect 4450 550 4460 570
rect 4160 540 4460 550
rect 4590 570 4890 580
rect 4590 550 4600 570
rect 4880 550 4890 570
rect 4590 540 4890 550
rect 50 440 1850 450
rect 50 420 410 440
rect 650 420 1850 440
rect 400 410 660 420
rect 60 380 360 390
rect 60 360 70 380
rect 350 360 660 380
rect 60 350 660 360
rect 60 280 660 310
rect 5060 430 5140 440
rect 5060 410 5070 430
rect 5130 410 5140 430
rect 5060 400 5140 410
rect 5060 350 5140 360
rect 3670 300 3970 340
rect 4160 300 4460 340
rect 4590 330 4890 340
rect 4590 310 4600 330
rect 4880 310 4890 330
rect 5060 330 5070 350
rect 5130 330 5140 350
rect 5060 320 5140 330
rect 4590 300 4890 310
rect 60 240 70 280
rect 40 230 70 240
rect 350 240 690 280
rect 350 230 1840 240
rect 40 210 1840 230
rect 40 100 1840 110
rect 40 70 50 100
rect 1820 70 1840 100
rect 40 60 1840 70
rect 3670 90 3970 100
rect 3670 70 3680 90
rect 3960 70 3970 90
rect 3670 60 3970 70
rect 4160 90 4460 100
rect 4160 70 4170 90
rect 4450 70 4460 90
rect 4160 60 4460 70
rect 4590 90 4890 100
rect 4590 70 4600 90
rect 4880 70 4890 90
rect 4590 60 4890 70
<< ndiffc >>
rect 2080 550 2360 570
rect 2880 550 3160 570
rect 5300 560 5580 580
rect 2080 310 2360 330
rect 2880 310 3160 330
rect 5300 310 5580 340
rect 5020 190 5080 210
rect 5020 110 5080 130
rect 2080 70 2660 90
rect 2880 70 3460 90
rect 5300 70 5580 90
<< pdiffc >>
rect 60 560 1840 580
rect 3680 550 3960 570
rect 4170 550 4450 570
rect 4600 550 4880 570
rect 410 420 650 440
rect 70 360 350 380
rect 5070 410 5130 430
rect 4600 310 4880 330
rect 5070 330 5130 350
rect 70 230 350 280
rect 50 70 1820 100
rect 3680 70 3960 90
rect 4170 70 4450 90
rect 4600 70 4880 90
<< psubdiff >>
rect 3290 500 3440 520
rect 3290 420 3310 500
rect 3420 420 3440 500
rect 3290 400 3440 420
rect 5660 500 5770 520
rect 5660 400 5680 500
rect 5750 400 5770 500
rect 5660 380 5770 400
<< nsubdiff >>
rect 5040 570 5180 590
rect 1100 360 1390 380
rect 1100 300 1120 360
rect 1370 300 1390 360
rect 5040 520 5060 570
rect 5160 520 5180 570
rect 5040 500 5180 520
rect 1100 280 1390 300
<< psubdiffcont >>
rect 3310 420 3420 500
rect 5680 400 5750 500
<< nsubdiffcont >>
rect 1120 300 1370 360
rect 5060 520 5160 570
<< poly >>
rect -40 540 50 550
rect -40 460 -30 540
rect 10 460 50 540
rect -40 450 50 460
rect 1850 450 1880 550
rect -30 340 60 350
rect -30 320 -20 340
rect 30 320 60 340
rect -30 310 60 320
rect 660 310 690 350
rect 2040 340 2070 540
rect 2370 510 2870 540
rect 2370 370 2440 510
rect 2800 370 2870 510
rect 2370 340 2870 370
rect 3170 340 3200 540
rect 3640 340 3670 540
rect 3970 480 4160 540
rect 3970 400 4020 480
rect 4100 400 4160 480
rect 3970 340 4160 400
rect 4460 340 4490 540
rect 4560 340 4590 540
rect 4890 510 4980 540
rect 4890 370 4920 510
rect 4970 370 4980 510
rect 5230 530 5290 550
rect 5160 460 5200 470
rect 5160 410 5170 460
rect 5190 410 5200 460
rect 5160 400 5200 410
rect 4890 340 4980 370
rect 5030 360 5060 400
rect 5140 360 5200 400
rect 5230 370 5240 530
rect 5270 370 5290 530
rect 5230 350 5290 370
rect 5590 350 5630 550
rect -40 200 40 210
rect -40 120 -30 200
rect 0 120 40 200
rect -40 110 40 120
rect 1840 110 1870 210
rect 2040 100 2070 300
rect 2670 260 2870 300
rect 2670 140 2720 260
rect 2820 140 2870 260
rect 2670 100 2870 140
rect 3470 100 3500 300
rect 3640 100 3670 300
rect 3970 100 4160 300
rect 4460 270 4590 300
rect 4460 130 4490 270
rect 4560 130 4590 270
rect 4460 100 4590 130
rect 4890 260 4960 300
rect 4890 130 4920 260
rect 4950 130 4960 260
rect 4990 140 5010 180
rect 5090 170 5190 180
rect 5090 150 5120 170
rect 5180 150 5190 170
rect 5090 140 5190 150
rect 4890 100 4960 130
rect 5250 100 5290 300
rect 5590 270 5680 300
rect 5590 130 5610 270
rect 5660 130 5680 270
rect 5590 100 5680 130
<< polycont >>
rect -30 460 10 540
rect -20 320 30 340
rect 2440 370 2800 510
rect 4020 400 4100 480
rect 4920 370 4970 510
rect 5170 410 5190 460
rect 5240 370 5270 530
rect -30 120 0 200
rect 2720 140 2820 260
rect 4490 130 4560 270
rect 4920 130 4950 260
rect 5120 150 5180 170
rect 5610 130 5660 270
<< locali >>
rect 50 580 1850 590
rect 5220 580 5590 590
rect 50 560 60 580
rect 1840 560 1850 580
rect 50 550 1850 560
rect 2070 570 2370 580
rect 2070 550 2080 570
rect 2360 550 2370 570
rect -40 540 20 550
rect 2070 540 2370 550
rect 2870 570 3610 580
rect 2870 550 2880 570
rect 3160 550 3610 570
rect 2870 540 3610 550
rect 3670 570 3970 580
rect 3670 550 3680 570
rect 3960 550 3970 570
rect 3670 540 3970 550
rect 4160 570 4460 580
rect 4160 550 4170 570
rect 4450 550 4460 570
rect 4160 540 4460 550
rect 4590 570 4890 580
rect 4590 550 4600 570
rect 4880 550 4890 570
rect 4590 540 4890 550
rect 5050 570 5170 580
rect -40 460 -30 540
rect 10 460 20 540
rect 3560 520 3610 540
rect 5050 520 5060 570
rect 5160 520 5170 570
rect -40 450 20 460
rect 2430 510 2810 520
rect 400 440 660 450
rect 400 420 410 440
rect 650 420 660 440
rect 60 400 110 410
rect 60 360 70 400
rect 100 390 110 400
rect 100 380 360 390
rect 350 360 360 380
rect 60 350 360 360
rect -30 340 40 350
rect -30 320 -20 340
rect 30 320 40 340
rect -30 310 40 320
rect 400 290 660 420
rect 2430 370 2440 510
rect 2800 370 2810 510
rect 1110 360 1380 370
rect 2430 360 2810 370
rect 3290 500 3440 520
rect 3290 420 3310 500
rect 3420 420 3440 500
rect 3290 390 3440 420
rect 3290 360 3340 390
rect 3390 360 3440 390
rect 1110 300 1120 360
rect 1370 300 1380 360
rect 3290 350 3440 360
rect 3560 480 4140 520
rect 3560 400 4020 480
rect 4100 400 4140 480
rect 3560 360 4140 400
rect 4910 510 4980 520
rect 5050 510 5170 520
rect 5220 560 5300 580
rect 5580 560 5590 580
rect 5220 550 5590 560
rect 5220 530 5290 550
rect 4910 370 4920 510
rect 4970 370 4980 510
rect 5160 460 5200 470
rect 5060 430 5140 440
rect 5060 410 5070 430
rect 5130 410 5140 430
rect 5060 400 5140 410
rect 5160 410 5170 460
rect 5190 410 5200 460
rect 5160 400 5200 410
rect 1110 290 1380 300
rect 1960 330 2380 340
rect 1960 310 2080 330
rect 2360 310 2380 330
rect 1960 300 2380 310
rect 2870 330 3170 340
rect 2870 310 2880 330
rect 3160 310 3170 330
rect 2870 300 3170 310
rect 60 280 660 290
rect 60 230 70 280
rect 350 230 660 280
rect 60 220 660 230
rect -40 200 10 210
rect -40 120 -30 200
rect 0 120 10 200
rect -40 110 10 120
rect 1960 110 2000 300
rect 2710 260 2830 270
rect 2710 140 2720 260
rect 2820 140 2830 260
rect 2710 130 2830 140
rect 40 100 2000 110
rect 3560 100 3610 360
rect 4910 340 4980 370
rect 5220 370 5240 530
rect 5270 370 5290 530
rect 5670 500 5760 510
rect 5670 400 5680 500
rect 5750 400 5760 500
rect 5670 390 5760 400
rect 5220 360 5270 370
rect 4590 330 4980 340
rect 4590 310 4600 330
rect 4880 310 4980 330
rect 5060 350 5270 360
rect 5060 330 5070 350
rect 5130 330 5270 350
rect 5060 320 5270 330
rect 5290 340 5590 350
rect 4590 300 4980 310
rect 5290 310 5300 340
rect 5580 310 5670 340
rect 5290 300 5670 310
rect 4480 270 4570 280
rect 5600 270 5670 300
rect 4480 130 4490 270
rect 4560 130 4570 270
rect 4480 100 4570 130
rect 4910 260 4960 270
rect 4910 130 4920 260
rect 4950 220 4960 260
rect 4950 210 5090 220
rect 4950 190 5020 210
rect 5080 190 5090 210
rect 4950 180 5090 190
rect 4950 130 4960 180
rect 5110 170 5190 180
rect 5110 150 5120 170
rect 5180 150 5190 170
rect 5110 140 5190 150
rect 4910 120 4960 130
rect 5010 130 5090 140
rect 5010 110 5020 130
rect 5080 110 5090 130
rect 5600 130 5610 270
rect 5660 130 5670 270
rect 5600 120 5670 130
rect 5010 100 5090 110
rect 40 70 50 100
rect 1820 70 2000 100
rect 40 60 2000 70
rect 2070 90 2670 100
rect 2070 70 2080 90
rect 2660 70 2670 90
rect 2070 60 2670 70
rect 2870 90 3470 100
rect 2870 70 2880 90
rect 3460 70 3470 90
rect 2870 60 3470 70
rect 3560 90 3970 100
rect 3560 70 3680 90
rect 3960 70 3970 90
rect 3560 60 3970 70
rect 4160 90 4460 100
rect 4160 70 4170 90
rect 4450 70 4460 90
rect 4160 60 4460 70
rect 4480 90 4890 100
rect 4480 70 4600 90
rect 4880 70 4890 90
rect 4480 60 4890 70
rect 5290 90 5590 100
rect 5290 70 5300 90
rect 5580 70 5590 90
rect 5290 60 5590 70
<< viali >>
rect 1800 560 1840 580
rect 2200 550 2250 570
rect 3800 550 3840 570
rect 4270 550 4310 570
rect 4710 550 4750 570
rect -30 470 10 520
rect 5090 520 5130 560
rect 70 380 100 400
rect 70 370 100 380
rect -20 320 10 340
rect 2570 410 2670 460
rect 3340 360 3390 390
rect 1230 300 1270 340
rect 5080 410 5120 430
rect 5170 420 5190 450
rect 2920 310 2960 330
rect -30 140 0 180
rect 2730 160 2810 240
rect 5700 420 5730 460
rect 5070 330 5130 350
rect 5140 150 5170 170
rect 5030 110 5070 130
rect 2270 70 2320 90
rect 3100 70 3150 90
rect 4260 70 4290 90
rect 5420 70 5470 90
<< metal1 >>
rect 1790 580 1850 590
rect 1790 550 1800 580
rect 1840 550 1850 580
rect -40 520 20 550
rect 1790 540 1850 550
rect 2190 550 2200 580
rect 2230 570 2260 580
rect 2250 550 2260 570
rect 2190 540 2260 550
rect 3790 550 3800 580
rect 3840 550 3850 580
rect 3790 540 3850 550
rect 4260 550 4270 580
rect 4310 550 4320 580
rect 4260 540 4320 550
rect 4700 550 4710 580
rect 4750 550 4760 580
rect 4700 540 4760 550
rect 5080 560 5140 570
rect -40 470 -30 520
rect 10 470 20 520
rect 5080 520 5090 560
rect 5130 520 5140 560
rect 5080 510 5140 520
rect -40 420 20 470
rect 2520 460 2740 490
rect 5690 460 5740 470
rect 2520 410 2570 460
rect 2670 420 4960 460
rect 5160 450 5200 460
rect 2670 410 2740 420
rect 60 400 110 410
rect 60 370 70 400
rect 100 370 110 400
rect 2520 390 2740 410
rect 3330 390 3400 400
rect 60 360 110 370
rect 3330 360 3340 390
rect 3390 360 3400 390
rect -30 340 20 360
rect 3330 350 3400 360
rect 4920 360 4960 420
rect 5070 410 5080 440
rect 5120 410 5130 440
rect 5160 420 5170 450
rect 5160 410 5200 420
rect 5690 420 5700 460
rect 5690 410 5740 420
rect 5070 400 5130 410
rect 4920 350 5140 360
rect -30 310 -20 340
rect 10 310 20 340
rect -30 300 20 310
rect 1220 340 1280 350
rect 1220 300 1230 340
rect 1270 300 1280 340
rect 2910 310 2920 340
rect 2960 310 2970 340
rect 4920 330 5070 350
rect 5130 330 5140 350
rect 4920 320 5140 330
rect 2910 300 2970 310
rect 1220 290 1280 300
rect 2720 240 2820 250
rect -40 180 10 240
rect -40 140 -30 180
rect 0 140 10 180
rect 2720 160 2730 240
rect 2810 160 2820 240
rect 2720 150 2820 160
rect 5130 150 5140 180
rect 5170 150 5180 180
rect 5130 140 5180 150
rect -40 110 10 140
rect 5020 130 5080 140
rect 4250 100 4310 110
rect 5020 100 5030 130
rect 5070 100 5080 130
rect 2260 90 2330 100
rect 2260 60 2270 90
rect 2320 70 2330 90
rect 2300 60 2330 70
rect 3090 90 3160 100
rect 3090 60 3100 90
rect 3150 70 3160 90
rect 3130 60 3160 70
rect 4250 70 4260 100
rect 4300 70 4310 100
rect 4250 60 4310 70
rect 5410 90 5480 100
rect 5410 60 5420 90
rect 5470 70 5480 90
rect 5460 60 5480 70
<< via1 >>
rect 1800 560 1840 580
rect 1800 550 1840 560
rect 2200 570 2230 580
rect 2200 550 2230 570
rect 3800 570 3840 580
rect 3800 550 3840 570
rect 4270 570 4310 580
rect 4270 550 4310 570
rect 4710 570 4750 580
rect 4710 550 4750 570
rect 5090 520 5130 560
rect 70 370 100 400
rect 3350 360 3380 390
rect 5080 430 5120 440
rect 5080 410 5120 430
rect 5170 420 5190 450
rect 5190 420 5200 450
rect 5700 420 5730 460
rect 5730 420 5740 460
rect -20 320 10 340
rect -20 310 10 320
rect 1230 300 1270 340
rect 2920 330 2960 340
rect 2920 310 2960 330
rect 2730 160 2810 240
rect 5140 170 5170 180
rect 5140 150 5170 170
rect 5030 110 5070 130
rect 5030 100 5070 110
rect 2270 70 2300 90
rect 2270 60 2300 70
rect 3100 70 3130 90
rect 3100 60 3130 70
rect 4260 90 4300 100
rect 4260 70 4290 90
rect 4290 70 4300 90
rect 5420 70 5460 90
rect 5420 60 5460 70
<< metal2 >>
rect -40 610 5780 650
rect 60 400 100 610
rect 60 370 70 400
rect 60 350 100 370
rect -30 340 20 350
rect 1220 340 1280 610
rect 3790 580 3850 610
rect -30 300 -20 340
rect 20 300 30 340
rect -20 290 30 300
rect 1220 300 1230 340
rect 1270 300 1280 340
rect 1790 550 1800 580
rect 1840 550 1850 580
rect 1790 340 1850 550
rect 2190 550 2200 580
rect 2230 550 2740 580
rect 2770 550 3610 580
rect 2190 540 3610 550
rect 3790 550 3800 580
rect 3840 550 3850 580
rect 4260 580 4320 610
rect 4260 550 4270 580
rect 4310 550 4320 580
rect 4700 580 4760 610
rect 4700 550 4710 580
rect 4750 550 4760 580
rect 3790 540 3850 550
rect 4700 540 4760 550
rect 5080 560 5140 610
rect 3340 390 3390 400
rect 3340 360 3350 390
rect 3380 360 3390 390
rect 1790 310 2920 340
rect 2960 310 2990 340
rect 1790 300 2990 310
rect 1220 290 1280 300
rect 2720 240 2820 250
rect 2720 160 2730 240
rect 2810 160 2820 240
rect 2720 150 2820 160
rect 2260 60 2270 90
rect 2300 60 2310 90
rect 2260 40 2310 60
rect 3090 60 3100 90
rect 3130 60 3140 90
rect 3090 40 3140 60
rect 3340 40 3390 360
rect 3560 100 3610 540
rect 5080 520 5090 560
rect 5130 520 5140 560
rect 5080 440 5140 520
rect 5120 410 5140 440
rect 5080 400 5140 410
rect 5160 460 5200 470
rect 5160 400 5200 420
rect 5690 460 5750 470
rect 5690 420 5700 460
rect 5740 420 5750 460
rect 5130 190 5190 200
rect 5130 150 5140 190
rect 5180 150 5190 190
rect 5130 140 5190 150
rect 5020 130 5080 140
rect 5020 100 5030 130
rect 5070 100 5080 130
rect 3560 70 4260 100
rect 4300 70 4460 100
rect 3560 60 4460 70
rect 5020 40 5080 100
rect 5410 60 5420 90
rect 5460 60 5470 90
rect 5410 40 5470 60
rect 5690 40 5750 420
rect -40 0 5780 40
<< via2 >>
rect -20 310 10 340
rect 10 310 20 340
rect -20 300 20 310
rect 2740 550 2770 580
rect 2730 160 2810 240
rect 5160 450 5200 460
rect 5160 420 5170 450
rect 5170 420 5200 450
rect 5140 180 5180 190
rect 5140 150 5170 180
rect 5170 150 5180 180
<< metal3 >>
rect 2730 580 5780 590
rect 2730 550 2740 580
rect 2770 550 5780 580
rect 2730 540 5780 550
rect 5150 460 5210 470
rect 5150 420 5160 460
rect 5200 420 5210 460
rect 5150 350 5210 420
rect -30 340 5230 350
rect -30 300 -20 340
rect 20 300 5230 340
rect -30 290 30 300
rect 2720 240 2820 250
rect 2720 160 2730 240
rect 2810 160 2820 240
rect 2720 150 2820 160
rect 5130 190 5190 200
rect 5130 150 5140 190
rect 5180 150 5190 190
rect 2750 70 2790 150
rect 5130 70 5190 150
rect 2750 40 5780 70
<< labels >>
rlabel metal1 -40 420 20 440 1 vin1
port 1 n
rlabel metal1 -40 220 10 240 1 vin2
port 2 n
rlabel metal1 -30 350 20 360 1 pbias
port 3 n
rlabel metal2 -40 610 -10 650 1 vdd
port 4 n
rlabel metal2 -40 0 -10 40 1 gnd
port 5 n
rlabel locali 400 320 660 370 1 nint
rlabel metal2 1880 300 1950 340 1 n14
rlabel locali 1960 160 2000 240 1 n23
rlabel locali 3290 540 3460 580 1 n810
rlabel pdiff 3670 300 3970 340 1 n68
rlabel pdiff 4160 300 4460 340 1 n57
rlabel pdiff 4590 300 4890 340 1 psc
rlabel poly 4890 100 4920 300 1 pcasc
rlabel ndiff 5290 300 5590 350 1 nsc
rlabel locali 5200 320 5270 360 1 ncasc
rlabel metal3 5760 40 5780 70 1 nbias
port 6 n
rlabel metal3 5750 540 5780 590 1 vout
port 7 n
<< end >>
