magic
tech sky130A
magscale 1 2
timestamp 1699666064
<< nwell >>
rect 200 -190 1910 310
rect 3180 -40 3900 760
<< nmos >>
rect 340 560 420 660
rect 1200 520 1300 760
rect 2480 40 2560 540
<< pmos >>
rect 450 40 1650 130
rect 3490 80 3580 580
<< ndiff >>
rect 270 630 340 660
rect 270 590 280 630
rect 320 590 340 630
rect 270 560 340 590
rect 420 630 490 660
rect 420 590 440 630
rect 480 590 490 630
rect 420 560 490 590
rect 1120 630 1200 760
rect 1120 580 1130 630
rect 1180 580 1200 630
rect 1120 520 1200 580
rect 1300 520 1380 760
rect 2410 230 2480 540
rect 2410 180 2420 230
rect 2460 180 2480 230
rect 2410 40 2480 180
rect 2560 230 2630 540
rect 2560 180 2580 230
rect 2620 180 2630 230
rect 2560 40 2630 180
<< pdiff >>
rect 330 110 450 130
rect 330 60 350 110
rect 410 60 450 110
rect 330 40 450 60
rect 1650 110 1770 130
rect 1650 60 1690 110
rect 1750 60 1770 110
rect 1650 40 1770 60
rect 3400 320 3490 580
rect 3400 210 3420 320
rect 3470 210 3490 320
rect 3400 80 3490 210
rect 3580 320 3670 580
rect 3580 210 3600 320
rect 3650 210 3670 320
rect 3580 80 3670 210
<< ndiffc >>
rect 280 590 320 630
rect 440 590 480 630
rect 1130 580 1180 630
rect 2420 180 2460 230
rect 2580 180 2620 230
<< pdiffc >>
rect 350 60 410 110
rect 1690 60 1750 110
rect 3420 210 3470 320
rect 3600 210 3650 320
<< psubdiff >>
rect 330 480 430 500
rect 330 440 360 480
rect 400 440 430 480
rect 330 420 430 440
rect 2480 -110 2580 -90
rect 2480 -150 2510 -110
rect 2550 -150 2580 -110
rect 2480 -170 2580 -150
<< nsubdiff >>
rect 3490 700 3610 720
rect 3490 660 3520 700
rect 3570 660 3610 700
rect 3490 640 3610 660
rect 240 260 1860 270
rect 240 220 930 260
rect 980 220 1860 260
rect 240 210 1860 220
rect 240 -90 270 210
rect 1830 -90 1860 210
rect 240 -150 1860 -90
<< psubdiffcont >>
rect 360 440 400 480
rect 2510 -150 2550 -110
<< nsubdiffcont >>
rect 3520 660 3570 700
rect 930 220 980 260
<< poly >>
rect 1200 840 1300 850
rect 1200 800 1230 840
rect 1270 800 1300 840
rect 1200 760 1300 800
rect 340 740 420 750
rect 340 700 360 740
rect 400 700 420 740
rect 340 660 420 700
rect 340 530 420 560
rect 2480 620 2560 630
rect 2480 580 2500 620
rect 2540 580 2560 620
rect 3490 580 3580 610
rect 2480 540 2560 580
rect 1200 490 1300 520
rect 450 130 1650 160
rect 450 10 1650 40
rect 910 -10 1010 10
rect 910 -50 940 -10
rect 980 -50 1010 -10
rect 910 -60 1010 -50
rect 2480 10 2560 40
rect 3490 30 3580 80
rect 3490 -10 3510 30
rect 3550 -10 3580 30
rect 3490 -20 3580 -10
<< polycont >>
rect 1230 800 1270 840
rect 360 700 400 740
rect 2500 580 2540 620
rect 940 -50 980 -10
rect 3510 -10 3550 30
<< locali >>
rect 1200 840 1300 850
rect 1200 800 1230 840
rect 1270 800 1300 840
rect 340 740 420 750
rect 340 700 360 740
rect 400 700 420 740
rect 280 630 340 660
rect 320 590 340 630
rect 280 560 340 590
rect 420 630 480 660
rect 420 590 440 630
rect 420 560 480 590
rect 1120 630 1200 760
rect 1120 580 1130 630
rect 1180 580 1200 630
rect 1120 520 1200 580
rect 1300 630 1380 760
rect 3490 700 3610 720
rect 3490 660 3520 700
rect 3570 660 3610 700
rect 3490 640 3610 660
rect 1300 580 1320 630
rect 1370 580 1380 630
rect 2480 620 2560 630
rect 2480 580 2500 620
rect 2540 580 2560 620
rect 1300 520 1380 580
rect 330 480 430 500
rect 330 440 360 480
rect 400 440 430 480
rect 330 420 430 440
rect 900 260 1020 270
rect 900 220 930 260
rect 980 220 1020 260
rect 900 210 1020 220
rect 2410 230 2480 540
rect 2410 180 2420 230
rect 2460 180 2480 230
rect 330 110 450 130
rect 330 60 350 110
rect 410 60 450 110
rect 330 40 450 60
rect 1650 110 1770 130
rect 1650 60 1690 110
rect 1750 60 1770 110
rect 1650 40 1770 60
rect 2410 40 2480 180
rect 2560 230 2630 540
rect 2560 180 2580 230
rect 2620 180 2630 230
rect 2560 40 2630 180
rect 3400 320 3490 580
rect 3400 210 3420 320
rect 3470 210 3490 320
rect 3400 80 3490 210
rect 3580 320 3670 580
rect 3580 210 3600 320
rect 3650 210 3670 320
rect 3580 80 3670 210
rect 3490 30 3580 40
rect 910 -10 1010 10
rect 910 -50 940 -10
rect 980 -50 1010 -10
rect 3490 -10 3510 30
rect 3550 -10 3580 30
rect 3490 -20 3580 -10
rect 910 -60 1010 -50
rect 2480 -110 2580 -90
rect 2480 -150 2510 -110
rect 2550 -150 2580 -110
rect 2480 -170 2580 -150
<< viali >>
rect 1230 800 1270 840
rect 360 700 400 740
rect 280 590 320 630
rect 440 590 480 630
rect 1130 580 1180 630
rect 3520 660 3570 700
rect 1320 580 1370 630
rect 2500 580 2540 620
rect 360 440 400 480
rect 930 220 980 260
rect 2420 180 2460 230
rect 350 60 410 110
rect 1690 60 1750 110
rect 2580 180 2620 230
rect 3420 210 3470 320
rect 3600 210 3650 320
rect 940 -50 980 -10
rect 3510 -10 3550 30
rect 2510 -150 2550 -110
<< metal1 >>
rect 200 960 4900 1000
rect 200 900 2100 960
rect 1200 840 1330 860
rect 1200 780 1230 840
rect 1300 780 1330 840
rect 1200 770 1330 780
rect 340 740 930 750
rect 340 700 360 740
rect 400 700 930 740
rect 340 690 930 700
rect 200 630 340 660
rect 200 590 280 630
rect 320 590 340 630
rect 200 560 340 590
rect 420 630 690 660
rect 420 590 440 630
rect 480 590 690 630
rect 420 560 690 590
rect 860 650 930 690
rect 1580 650 1650 900
rect 2000 890 2100 900
rect 2190 900 4900 960
rect 2190 890 2320 900
rect 2000 870 2320 890
rect 2720 800 2860 820
rect 2720 720 2740 800
rect 2840 720 2860 800
rect 3660 720 3770 900
rect 2720 700 2860 720
rect 3490 700 3770 720
rect 860 632 1200 650
rect 860 573 1111 632
rect 1181 573 1200 632
rect 860 560 1200 573
rect 1300 630 1650 650
rect 1300 580 1320 630
rect 1370 580 1650 630
rect 1300 560 1650 580
rect 2480 630 2600 640
rect 2480 570 2490 630
rect 2550 570 2600 630
rect 2480 560 2600 570
rect 200 500 290 560
rect 200 480 430 500
rect 200 440 360 480
rect 400 440 430 480
rect 200 420 430 440
rect 630 470 690 560
rect 200 -200 270 420
rect 630 380 2250 470
rect 900 260 1780 270
rect 900 220 930 260
rect 980 220 1780 260
rect 900 210 1780 220
rect 1690 130 1780 210
rect 2180 240 2250 380
rect 2740 240 2840 700
rect 3490 660 3520 700
rect 3570 660 3770 700
rect 3490 640 3770 660
rect 3660 340 3770 640
rect 3370 320 3490 340
rect 3370 240 3420 320
rect 2180 230 2480 240
rect 2180 180 2420 230
rect 2460 180 2480 230
rect 2180 160 2480 180
rect 2560 230 3420 240
rect 2560 180 2580 230
rect 2620 210 3420 230
rect 3470 210 3490 320
rect 2620 190 3490 210
rect 3580 320 3770 340
rect 3580 210 3600 320
rect 3650 210 3770 320
rect 3580 190 3770 210
rect 2620 180 3470 190
rect 2560 170 3470 180
rect 2560 160 2650 170
rect 330 110 450 130
rect 330 60 350 110
rect 410 60 450 110
rect 330 40 450 60
rect 1650 110 1780 130
rect 1650 60 1690 110
rect 1750 60 1780 110
rect 1650 40 1780 60
rect 330 10 440 40
rect 330 0 1010 10
rect 330 -60 930 0
rect 1000 -60 1010 0
rect 1690 -10 1780 40
rect 2740 -10 2800 170
rect 1690 -60 2800 -10
rect 3490 -20 3500 40
rect 3560 -20 3580 40
rect 2480 -110 2580 -90
rect 2480 -150 2510 -110
rect 2550 -150 2580 -110
rect 2480 -200 2580 -150
rect 200 -300 4900 -200
<< via1 >>
rect 1230 800 1270 840
rect 1270 800 1300 840
rect 1230 780 1300 800
rect 2100 890 2190 960
rect 2740 720 2840 800
rect 1111 630 1181 632
rect 1111 580 1130 630
rect 1130 580 1180 630
rect 1180 580 1181 630
rect 1111 573 1181 580
rect 2490 620 2550 630
rect 2490 580 2500 620
rect 2500 580 2540 620
rect 2540 580 2550 620
rect 2490 570 2550 580
rect 930 -10 1000 0
rect 930 -50 940 -10
rect 940 -50 980 -10
rect 980 -50 1000 -10
rect 930 -60 1000 -50
rect 3500 30 3560 40
rect 3500 -10 3510 30
rect 3510 -10 3550 30
rect 3550 -10 3560 30
rect 3500 -20 3560 -10
<< metal2 >>
rect 2090 990 2300 1000
rect 2090 960 2180 990
rect 2090 890 2100 960
rect 2250 930 2300 990
rect 2190 890 2300 930
rect 910 880 1330 890
rect 2090 880 2300 890
rect 2720 990 4740 1000
rect 2720 930 4600 990
rect 4680 930 4740 990
rect 910 820 1010 880
rect 1080 840 1330 880
rect 1080 820 1230 840
rect 910 780 1230 820
rect 1300 780 1330 840
rect 910 760 1330 780
rect 2720 870 4740 930
rect 2720 800 4900 870
rect 910 0 1020 760
rect 2720 720 2740 800
rect 2840 720 2860 800
rect 2720 700 2860 720
rect 1080 632 1193 650
rect 1080 573 1111 632
rect 1181 573 1193 632
rect 1080 464 1193 573
rect 2480 630 4900 640
rect 2480 570 2490 630
rect 2550 570 4900 630
rect 2480 560 4900 570
rect 1079 387 4900 464
rect 910 -60 930 0
rect 1000 -60 1020 0
rect 3490 40 4900 50
rect 3490 -20 3500 40
rect 3560 -20 4900 40
rect 910 -80 1020 -60
<< via2 >>
rect 2180 960 2250 990
rect 2180 930 2190 960
rect 2190 930 2250 960
rect 4600 930 4680 990
rect 1010 820 1080 880
<< metal3 >>
rect 2130 990 2300 1000
rect 2130 920 2180 990
rect 2260 920 2300 990
rect 4560 994 4710 1000
rect 4560 926 4598 994
rect 4682 926 4710 994
rect 4560 920 4710 926
rect 890 880 1370 900
rect 890 840 1010 880
rect 160 820 1010 840
rect 1080 840 1370 880
rect 1080 820 4840 840
rect 160 -240 4840 820
rect 4340 -260 4840 -240
<< via3 >>
rect 2180 930 2250 990
rect 2250 930 2260 990
rect 2180 920 2260 930
rect 4598 990 4682 994
rect 4598 930 4600 990
rect 4600 930 4680 990
rect 4680 930 4682 990
rect 4598 926 4682 930
<< mimcap >>
rect 200 120 4200 800
rect 200 -80 2060 120
rect 2280 -80 4200 120
rect 200 -200 4200 -80
rect 4380 120 4780 800
rect 4380 -100 4440 120
rect 4680 -100 4780 120
rect 4380 -200 4780 -100
<< mimcapcontact >>
rect 2060 -80 2280 120
rect 4440 -100 4680 120
<< metal4 >>
rect 2000 990 2320 1000
rect 2000 920 2180 990
rect 2260 920 2320 990
rect 4560 994 4710 1000
rect 4560 960 4598 994
rect 2000 120 2320 920
rect 2000 -80 2060 120
rect 2280 -80 2320 120
rect 2000 -300 2320 -80
rect 4400 926 4598 960
rect 4682 960 4710 994
rect 4682 926 4740 960
rect 4400 120 4740 926
rect 4400 -100 4440 120
rect 4680 -100 4740 120
rect 4400 -280 4740 -100
<< labels >>
rlabel metal1 4845 937 4845 937 1 VDD
rlabel metal1 4860 -266 4860 -266 1 GND
rlabel metal2 4886 836 4886 836 1 VOUT
rlabel metal2 4886 600 4887 601 1 VCASN
rlabel metal2 4875 423 4875 423 1 IN
rlabel metal2 4870 10 4870 10 1 PBIAS
<< end >>
