magic
tech sky130A
timestamp 1702481431
<< nwell >>
rect -13 639 5246 640
rect -13 471 5271 639
rect -13 208 5246 471
rect -13 160 2172 208
<< nmos >>
rect -654 449 -614 579
rect -584 449 -544 579
rect -514 449 -474 579
rect -444 449 -404 579
rect -374 449 -334 579
rect -185 470 -145 550
rect -553 153 -473 173
rect -259 76 -219 276
rect -189 76 -149 276
rect 155 45 215 120
rect 245 45 305 120
rect 335 45 395 120
rect 425 45 485 120
rect 515 45 575 120
rect 605 45 665 120
rect 695 45 755 120
rect 785 45 845 120
rect 1295 45 1355 120
rect 1385 45 1445 120
rect 1475 45 1535 120
rect 1565 45 1625 120
rect 1655 45 1715 120
rect 1745 45 1805 120
rect 1835 45 1895 120
rect 1925 45 1985 120
rect 2249 39 2309 164
rect 2339 39 2399 164
rect 2429 39 2489 164
rect 2519 39 2579 164
rect 2609 39 2669 164
rect 2699 39 2759 164
rect 2789 39 2849 164
rect 2879 39 2939 164
rect 2969 39 3029 164
rect 3059 39 3119 164
rect 3149 39 3209 164
rect 3239 39 3299 164
rect 3329 39 3389 164
rect 3419 39 3479 164
rect 3509 39 3569 164
rect 3599 39 3659 164
rect 3759 39 3819 164
rect 3849 39 3909 164
rect 3939 39 3999 164
rect 4029 39 4089 164
rect 4119 39 4179 164
rect 4209 39 4269 164
rect 4299 39 4359 164
rect 4389 39 4449 164
rect 4479 39 4539 164
rect 4569 39 4629 164
rect 4659 39 4719 164
rect 4749 39 4809 164
rect 4839 39 4899 164
rect 4929 39 4989 164
rect 5019 39 5079 164
rect 5109 39 5169 164
<< pmos >>
rect 70 441 110 591
rect 150 441 190 591
rect 230 441 270 591
rect 310 441 350 591
rect 390 441 430 591
rect 470 441 510 591
rect 550 441 590 591
rect 630 441 670 591
rect 710 441 750 591
rect 790 441 830 591
rect 870 441 910 591
rect 950 441 990 591
rect 1030 441 1070 591
rect 1110 441 1150 591
rect 1190 441 1230 591
rect 1270 441 1310 591
rect 1350 441 1390 591
rect 1430 441 1470 591
rect 1510 441 1550 591
rect 1590 441 1630 591
rect 1670 441 1710 591
rect 1750 441 1790 591
rect 1830 441 1870 591
rect 1910 441 1950 591
rect 1990 441 2030 591
rect 2070 441 2110 591
rect 2249 459 2309 584
rect 2339 459 2399 584
rect 2429 459 2489 584
rect 2519 459 2579 584
rect 2609 459 2669 584
rect 2699 459 2759 584
rect 2789 459 2849 584
rect 2879 459 2939 584
rect 2969 459 3029 584
rect 3059 459 3119 584
rect 3149 459 3209 584
rect 3239 459 3299 584
rect 3329 459 3389 584
rect 3419 459 3479 584
rect 3509 459 3569 584
rect 3599 459 3659 584
rect 3759 459 3819 584
rect 3849 459 3909 584
rect 3939 459 3999 584
rect 4029 459 4089 584
rect 4119 459 4179 584
rect 4209 459 4269 584
rect 4299 459 4359 584
rect 4389 459 4449 584
rect 4479 459 4539 584
rect 4569 459 4629 584
rect 4659 459 4719 584
rect 4749 459 4809 584
rect 4839 459 4899 584
rect 4929 459 4989 584
rect 5019 459 5079 584
rect 5109 459 5169 584
rect 51 205 71 355
rect 101 205 121 355
rect 151 205 171 355
rect 201 205 221 355
rect 251 205 271 355
rect 301 205 321 355
rect 351 205 371 355
rect 401 205 421 355
rect 451 205 471 355
rect 501 205 521 355
rect 551 205 571 355
rect 601 205 621 355
rect 651 205 671 355
rect 701 205 721 355
rect 751 205 771 355
rect 801 205 821 355
rect 851 205 871 355
rect 901 205 921 355
rect 951 205 971 355
rect 1001 205 1021 355
rect 1151 205 1171 355
rect 1201 205 1221 355
rect 1251 205 1271 355
rect 1301 205 1321 355
rect 1351 205 1371 355
rect 1401 205 1421 355
rect 1451 205 1471 355
rect 1501 205 1521 355
rect 1551 205 1571 355
rect 1601 205 1621 355
rect 1651 205 1671 355
rect 1701 205 1721 355
rect 1751 205 1771 355
rect 1801 205 1821 355
rect 1851 205 1871 355
rect 1901 205 1921 355
rect 1951 205 1971 355
rect 2001 205 2021 355
rect 2051 205 2071 355
rect 2101 205 2121 355
rect 2249 244 2309 369
rect 2339 244 2399 369
rect 2429 244 2489 369
rect 2519 244 2579 369
rect 2609 244 2669 369
rect 2699 244 2759 369
rect 2789 244 2849 369
rect 2879 244 2939 369
rect 2969 244 3029 369
rect 3059 244 3119 369
rect 3149 244 3209 369
rect 3239 244 3299 369
rect 3329 244 3389 369
rect 3419 244 3479 369
rect 3509 244 3569 369
rect 3599 244 3659 369
rect 3759 244 3819 369
rect 3849 244 3909 369
rect 3939 244 3999 369
rect 4029 244 4089 369
rect 4119 244 4179 369
rect 4209 244 4269 369
rect 4299 244 4359 369
rect 4389 244 4449 369
rect 4479 244 4539 369
rect 4569 244 4629 369
rect 4659 244 4719 369
rect 4749 244 4809 369
rect 4839 244 4899 369
rect 4929 244 4989 369
rect 5019 244 5079 369
rect 5109 244 5169 369
<< ndiff >>
rect -684 563 -654 579
rect -684 463 -677 563
rect -660 463 -654 563
rect -684 449 -654 463
rect -614 563 -584 579
rect -614 463 -607 563
rect -590 463 -584 563
rect -614 449 -584 463
rect -544 563 -514 579
rect -544 463 -537 563
rect -520 463 -514 563
rect -544 449 -514 463
rect -474 563 -444 579
rect -474 463 -467 563
rect -450 463 -444 563
rect -474 449 -444 463
rect -404 563 -374 579
rect -404 463 -397 563
rect -380 463 -374 563
rect -404 449 -374 463
rect -334 563 -304 579
rect -334 463 -327 563
rect -310 463 -304 563
rect -215 542 -185 550
rect -215 478 -209 542
rect -191 478 -185 542
rect -215 470 -185 478
rect -145 542 -115 550
rect -145 478 -139 542
rect -121 478 -115 542
rect -145 470 -115 478
rect -334 449 -304 463
rect -289 261 -259 276
rect -613 196 -583 214
rect -613 130 -607 196
rect -589 173 -583 196
rect -443 196 -413 214
rect -443 173 -437 196
rect -589 153 -553 173
rect -473 153 -437 173
rect -589 130 -583 153
rect -613 114 -583 130
rect -443 130 -437 153
rect -419 130 -413 196
rect -443 114 -413 130
rect -289 92 -282 261
rect -265 92 -259 261
rect -289 76 -259 92
rect -219 261 -189 276
rect -219 92 -212 261
rect -195 92 -189 261
rect -219 76 -189 92
rect -149 261 -119 276
rect -149 92 -142 261
rect -125 92 -119 261
rect 2219 151 2249 164
rect -149 76 -119 92
rect 125 106 155 120
rect 125 58 131 106
rect 149 58 155 106
rect 125 45 155 58
rect 215 106 245 120
rect 215 58 221 106
rect 239 58 245 106
rect 215 45 245 58
rect 305 106 335 120
rect 305 58 311 106
rect 329 58 335 106
rect 305 45 335 58
rect 395 106 425 120
rect 395 58 401 106
rect 419 58 425 106
rect 395 45 425 58
rect 485 106 515 120
rect 485 58 491 106
rect 509 58 515 106
rect 485 45 515 58
rect 575 106 605 120
rect 575 58 581 106
rect 599 58 605 106
rect 575 45 605 58
rect 665 106 695 120
rect 665 58 671 106
rect 689 58 695 106
rect 665 45 695 58
rect 755 106 785 120
rect 755 58 761 106
rect 779 58 785 106
rect 755 45 785 58
rect 845 106 875 120
rect 845 58 851 106
rect 869 58 875 106
rect 845 45 875 58
rect 1265 106 1295 120
rect 1265 58 1271 106
rect 1289 58 1295 106
rect 1265 45 1295 58
rect 1355 106 1385 120
rect 1355 58 1361 106
rect 1379 58 1385 106
rect 1355 45 1385 58
rect 1445 106 1475 120
rect 1445 58 1451 106
rect 1469 58 1475 106
rect 1445 45 1475 58
rect 1535 106 1565 120
rect 1535 58 1541 106
rect 1559 58 1565 106
rect 1535 45 1565 58
rect 1625 106 1655 120
rect 1625 58 1631 106
rect 1649 58 1655 106
rect 1625 45 1655 58
rect 1715 106 1745 120
rect 1715 58 1721 106
rect 1739 58 1745 106
rect 1715 45 1745 58
rect 1805 106 1835 120
rect 1805 58 1811 106
rect 1829 58 1835 106
rect 1805 45 1835 58
rect 1895 106 1925 120
rect 1895 58 1901 106
rect 1919 58 1925 106
rect 1895 45 1925 58
rect 1985 106 2015 120
rect 1985 58 1991 106
rect 2009 58 2015 106
rect 1985 45 2015 58
rect 2219 51 2225 151
rect 2243 51 2249 151
rect 2219 39 2249 51
rect 2309 151 2339 164
rect 2309 51 2315 151
rect 2333 51 2339 151
rect 2309 39 2339 51
rect 2399 151 2429 164
rect 2399 51 2405 151
rect 2423 51 2429 151
rect 2399 39 2429 51
rect 2489 151 2519 164
rect 2489 51 2495 151
rect 2513 51 2519 151
rect 2489 39 2519 51
rect 2579 151 2609 164
rect 2579 51 2585 151
rect 2603 51 2609 151
rect 2579 39 2609 51
rect 2669 151 2699 164
rect 2669 51 2675 151
rect 2693 51 2699 151
rect 2669 39 2699 51
rect 2759 151 2789 164
rect 2759 51 2765 151
rect 2783 51 2789 151
rect 2759 39 2789 51
rect 2849 151 2879 164
rect 2849 51 2855 151
rect 2873 51 2879 151
rect 2849 39 2879 51
rect 2939 151 2969 164
rect 2939 51 2945 151
rect 2963 51 2969 151
rect 2939 39 2969 51
rect 3029 151 3059 164
rect 3029 51 3035 151
rect 3053 51 3059 151
rect 3029 39 3059 51
rect 3119 151 3149 164
rect 3119 51 3125 151
rect 3143 51 3149 151
rect 3119 39 3149 51
rect 3209 151 3239 164
rect 3209 51 3215 151
rect 3233 51 3239 151
rect 3209 39 3239 51
rect 3299 151 3329 164
rect 3299 51 3305 151
rect 3323 51 3329 151
rect 3299 39 3329 51
rect 3389 151 3419 164
rect 3389 51 3395 151
rect 3413 51 3419 151
rect 3389 39 3419 51
rect 3479 151 3509 164
rect 3479 51 3485 151
rect 3503 51 3509 151
rect 3479 39 3509 51
rect 3569 151 3599 164
rect 3569 51 3575 151
rect 3593 51 3599 151
rect 3569 39 3599 51
rect 3659 151 3689 164
rect 3659 51 3665 151
rect 3683 51 3689 151
rect 3659 39 3689 51
rect 3729 151 3759 164
rect 3729 51 3735 151
rect 3753 51 3759 151
rect 3729 39 3759 51
rect 3819 151 3849 164
rect 3819 51 3825 151
rect 3843 51 3849 151
rect 3819 39 3849 51
rect 3909 151 3939 164
rect 3909 51 3915 151
rect 3933 51 3939 151
rect 3909 39 3939 51
rect 3999 151 4029 164
rect 3999 51 4005 151
rect 4023 51 4029 151
rect 3999 39 4029 51
rect 4089 151 4119 164
rect 4089 51 4095 151
rect 4113 51 4119 151
rect 4089 39 4119 51
rect 4179 151 4209 164
rect 4179 51 4185 151
rect 4203 51 4209 151
rect 4179 39 4209 51
rect 4269 151 4299 164
rect 4269 51 4275 151
rect 4293 51 4299 151
rect 4269 39 4299 51
rect 4359 151 4389 164
rect 4359 51 4365 151
rect 4383 51 4389 151
rect 4359 39 4389 51
rect 4449 151 4479 164
rect 4449 51 4455 151
rect 4473 51 4479 151
rect 4449 39 4479 51
rect 4539 151 4569 164
rect 4539 51 4545 151
rect 4563 51 4569 151
rect 4539 39 4569 51
rect 4629 151 4659 164
rect 4629 51 4635 151
rect 4653 51 4659 151
rect 4629 39 4659 51
rect 4719 151 4749 164
rect 4719 51 4725 151
rect 4743 51 4749 151
rect 4719 39 4749 51
rect 4809 151 4839 164
rect 4809 51 4815 151
rect 4833 51 4839 151
rect 4809 39 4839 51
rect 4899 151 4929 164
rect 4899 51 4905 151
rect 4923 51 4929 151
rect 4899 39 4929 51
rect 4989 151 5019 164
rect 4989 51 4995 151
rect 5013 51 5019 151
rect 4989 39 5019 51
rect 5079 151 5109 164
rect 5079 51 5085 151
rect 5103 51 5109 151
rect 5079 39 5109 51
rect 5169 151 5199 164
rect 5169 51 5175 151
rect 5193 51 5199 151
rect 5169 39 5199 51
<< pdiff >>
rect 30 582 70 591
rect 30 449 40 582
rect 61 449 70 582
rect 30 441 70 449
rect 110 582 150 591
rect 110 449 120 582
rect 141 449 150 582
rect 110 441 150 449
rect 190 582 230 591
rect 190 449 200 582
rect 221 449 230 582
rect 190 441 230 449
rect 270 582 310 591
rect 270 449 280 582
rect 301 449 310 582
rect 270 441 310 449
rect 350 582 390 591
rect 350 449 360 582
rect 381 449 390 582
rect 350 441 390 449
rect 430 582 470 591
rect 430 449 440 582
rect 461 449 470 582
rect 430 441 470 449
rect 510 582 550 591
rect 510 449 520 582
rect 541 449 550 582
rect 510 441 550 449
rect 590 582 630 591
rect 590 449 600 582
rect 621 449 630 582
rect 590 441 630 449
rect 670 582 710 591
rect 670 449 680 582
rect 701 449 710 582
rect 670 441 710 449
rect 750 582 790 591
rect 750 449 760 582
rect 781 449 790 582
rect 750 441 790 449
rect 830 582 870 591
rect 830 449 840 582
rect 861 449 870 582
rect 830 441 870 449
rect 910 582 950 591
rect 910 449 920 582
rect 941 449 950 582
rect 910 441 950 449
rect 990 582 1030 591
rect 990 449 1000 582
rect 1021 449 1030 582
rect 990 441 1030 449
rect 1070 582 1110 591
rect 1070 449 1080 582
rect 1101 449 1110 582
rect 1070 441 1110 449
rect 1150 582 1190 591
rect 1150 449 1160 582
rect 1181 449 1190 582
rect 1150 441 1190 449
rect 1230 582 1270 591
rect 1230 449 1240 582
rect 1261 449 1270 582
rect 1230 441 1270 449
rect 1310 582 1350 591
rect 1310 449 1320 582
rect 1341 449 1350 582
rect 1310 441 1350 449
rect 1390 582 1430 591
rect 1390 449 1400 582
rect 1421 449 1430 582
rect 1390 441 1430 449
rect 1470 582 1510 591
rect 1470 449 1480 582
rect 1501 449 1510 582
rect 1470 441 1510 449
rect 1550 582 1590 591
rect 1550 449 1560 582
rect 1581 449 1590 582
rect 1550 441 1590 449
rect 1630 582 1670 591
rect 1630 449 1640 582
rect 1661 449 1670 582
rect 1630 441 1670 449
rect 1710 582 1750 591
rect 1710 449 1720 582
rect 1741 449 1750 582
rect 1710 441 1750 449
rect 1790 582 1830 591
rect 1790 449 1800 582
rect 1821 449 1830 582
rect 1790 441 1830 449
rect 1870 582 1910 591
rect 1870 449 1880 582
rect 1901 449 1910 582
rect 1870 441 1910 449
rect 1950 582 1990 591
rect 1950 449 1960 582
rect 1981 449 1990 582
rect 1950 441 1990 449
rect 2030 582 2070 591
rect 2030 449 2040 582
rect 2061 449 2070 582
rect 2030 441 2070 449
rect 2110 582 2150 591
rect 2110 449 2120 582
rect 2141 449 2150 582
rect 2219 571 2249 584
rect 2219 471 2225 571
rect 2243 471 2249 571
rect 2219 459 2249 471
rect 2309 571 2339 584
rect 2309 471 2315 571
rect 2333 471 2339 571
rect 2309 459 2339 471
rect 2399 571 2429 584
rect 2399 471 2405 571
rect 2423 471 2429 571
rect 2399 459 2429 471
rect 2489 571 2519 584
rect 2489 471 2495 571
rect 2513 471 2519 571
rect 2489 459 2519 471
rect 2579 571 2609 584
rect 2579 471 2585 571
rect 2603 471 2609 571
rect 2579 459 2609 471
rect 2669 571 2699 584
rect 2669 471 2675 571
rect 2693 471 2699 571
rect 2669 459 2699 471
rect 2759 571 2789 584
rect 2759 471 2765 571
rect 2783 471 2789 571
rect 2759 459 2789 471
rect 2849 571 2879 584
rect 2849 471 2855 571
rect 2873 471 2879 571
rect 2849 459 2879 471
rect 2939 571 2969 584
rect 2939 471 2945 571
rect 2963 471 2969 571
rect 2939 459 2969 471
rect 3029 571 3059 584
rect 3029 471 3035 571
rect 3053 471 3059 571
rect 3029 459 3059 471
rect 3119 571 3149 584
rect 3119 471 3125 571
rect 3143 471 3149 571
rect 3119 459 3149 471
rect 3209 571 3239 584
rect 3209 471 3215 571
rect 3233 471 3239 571
rect 3209 459 3239 471
rect 3299 571 3329 584
rect 3299 471 3305 571
rect 3323 471 3329 571
rect 3299 459 3329 471
rect 3389 571 3419 584
rect 3389 471 3395 571
rect 3413 471 3419 571
rect 3389 459 3419 471
rect 3479 571 3509 584
rect 3479 471 3485 571
rect 3503 471 3509 571
rect 3479 459 3509 471
rect 3569 571 3599 584
rect 3569 471 3575 571
rect 3593 471 3599 571
rect 3569 459 3599 471
rect 3659 571 3689 584
rect 3659 471 3665 571
rect 3683 471 3689 571
rect 3659 459 3689 471
rect 3729 571 3759 584
rect 3729 471 3735 571
rect 3753 471 3759 571
rect 3729 459 3759 471
rect 3819 571 3849 584
rect 3819 471 3825 571
rect 3843 471 3849 571
rect 3819 459 3849 471
rect 3909 571 3939 584
rect 3909 471 3915 571
rect 3933 471 3939 571
rect 3909 459 3939 471
rect 3999 571 4029 584
rect 3999 471 4005 571
rect 4023 471 4029 571
rect 3999 459 4029 471
rect 4089 571 4119 584
rect 4089 471 4095 571
rect 4113 471 4119 571
rect 4089 459 4119 471
rect 4179 571 4209 584
rect 4179 471 4185 571
rect 4203 471 4209 571
rect 4179 459 4209 471
rect 4269 571 4299 584
rect 4269 471 4275 571
rect 4293 471 4299 571
rect 4269 459 4299 471
rect 4359 571 4389 584
rect 4359 471 4365 571
rect 4383 471 4389 571
rect 4359 459 4389 471
rect 4449 571 4479 584
rect 4449 471 4455 571
rect 4473 471 4479 571
rect 4449 459 4479 471
rect 4539 571 4569 584
rect 4539 471 4545 571
rect 4563 471 4569 571
rect 4539 459 4569 471
rect 4629 571 4659 584
rect 4629 471 4635 571
rect 4653 471 4659 571
rect 4629 459 4659 471
rect 4719 571 4749 584
rect 4719 471 4725 571
rect 4743 471 4749 571
rect 4719 459 4749 471
rect 4809 571 4839 584
rect 4809 471 4815 571
rect 4833 471 4839 571
rect 4809 459 4839 471
rect 4899 571 4929 584
rect 4899 471 4905 571
rect 4923 471 4929 571
rect 4899 459 4929 471
rect 4989 571 5019 584
rect 4989 471 4995 571
rect 5013 471 5019 571
rect 4989 459 5019 471
rect 5079 571 5109 584
rect 5079 471 5085 571
rect 5103 471 5109 571
rect 5079 459 5109 471
rect 5169 571 5199 584
rect 5169 471 5175 571
rect 5193 471 5199 571
rect 5169 459 5199 471
rect 2110 441 2150 449
rect 2219 356 2249 369
rect 21 335 51 355
rect 21 226 28 335
rect 45 226 51 335
rect 21 205 51 226
rect 71 335 101 355
rect 71 226 78 335
rect 95 226 101 335
rect 71 205 101 226
rect 121 335 151 355
rect 121 226 128 335
rect 145 226 151 335
rect 121 205 151 226
rect 171 335 201 355
rect 171 226 178 335
rect 195 226 201 335
rect 171 205 201 226
rect 221 335 251 355
rect 221 226 228 335
rect 245 226 251 335
rect 221 205 251 226
rect 271 335 301 355
rect 271 226 278 335
rect 295 226 301 335
rect 271 205 301 226
rect 321 335 351 355
rect 321 226 328 335
rect 345 226 351 335
rect 321 205 351 226
rect 371 335 401 355
rect 371 226 378 335
rect 395 226 401 335
rect 371 205 401 226
rect 421 335 451 355
rect 421 226 428 335
rect 445 226 451 335
rect 421 205 451 226
rect 471 335 501 355
rect 471 226 478 335
rect 495 226 501 335
rect 471 205 501 226
rect 521 335 551 355
rect 521 226 528 335
rect 545 226 551 335
rect 521 205 551 226
rect 571 335 601 355
rect 571 226 578 335
rect 595 226 601 335
rect 571 205 601 226
rect 621 335 651 355
rect 621 226 628 335
rect 645 226 651 335
rect 621 205 651 226
rect 671 335 701 355
rect 671 226 678 335
rect 695 226 701 335
rect 671 205 701 226
rect 721 335 751 355
rect 721 226 728 335
rect 745 226 751 335
rect 721 205 751 226
rect 771 335 801 355
rect 771 226 778 335
rect 795 226 801 335
rect 771 205 801 226
rect 821 335 851 355
rect 821 226 828 335
rect 845 226 851 335
rect 821 205 851 226
rect 871 335 901 355
rect 871 226 878 335
rect 895 226 901 335
rect 871 205 901 226
rect 921 335 951 355
rect 921 226 928 335
rect 945 226 951 335
rect 921 205 951 226
rect 971 335 1001 355
rect 971 226 978 335
rect 995 226 1001 335
rect 971 205 1001 226
rect 1021 335 1051 355
rect 1021 226 1028 335
rect 1045 226 1051 335
rect 1021 205 1051 226
rect 1121 335 1151 355
rect 1121 226 1128 335
rect 1145 226 1151 335
rect 1121 205 1151 226
rect 1171 335 1201 355
rect 1171 226 1178 335
rect 1195 226 1201 335
rect 1171 205 1201 226
rect 1221 335 1251 355
rect 1221 226 1228 335
rect 1245 226 1251 335
rect 1221 205 1251 226
rect 1271 335 1301 355
rect 1271 226 1278 335
rect 1295 226 1301 335
rect 1271 205 1301 226
rect 1321 335 1351 355
rect 1321 226 1328 335
rect 1345 226 1351 335
rect 1321 205 1351 226
rect 1371 335 1401 355
rect 1371 226 1378 335
rect 1395 226 1401 335
rect 1371 205 1401 226
rect 1421 335 1451 355
rect 1421 226 1428 335
rect 1445 226 1451 335
rect 1421 205 1451 226
rect 1471 335 1501 355
rect 1471 226 1478 335
rect 1495 226 1501 335
rect 1471 205 1501 226
rect 1521 335 1551 355
rect 1521 226 1528 335
rect 1545 226 1551 335
rect 1521 205 1551 226
rect 1571 335 1601 355
rect 1571 226 1578 335
rect 1595 226 1601 335
rect 1571 205 1601 226
rect 1621 335 1651 355
rect 1621 226 1628 335
rect 1645 226 1651 335
rect 1621 205 1651 226
rect 1671 335 1701 355
rect 1671 226 1678 335
rect 1695 226 1701 335
rect 1671 205 1701 226
rect 1721 335 1751 355
rect 1721 226 1728 335
rect 1745 226 1751 335
rect 1721 205 1751 226
rect 1771 335 1801 355
rect 1771 226 1778 335
rect 1795 226 1801 335
rect 1771 205 1801 226
rect 1821 335 1851 355
rect 1821 226 1828 335
rect 1845 226 1851 335
rect 1821 205 1851 226
rect 1871 335 1901 355
rect 1871 226 1878 335
rect 1895 226 1901 335
rect 1871 205 1901 226
rect 1921 335 1951 355
rect 1921 226 1928 335
rect 1945 226 1951 335
rect 1921 205 1951 226
rect 1971 335 2001 355
rect 1971 226 1978 335
rect 1995 226 2001 335
rect 1971 205 2001 226
rect 2021 335 2051 355
rect 2021 226 2028 335
rect 2045 226 2051 335
rect 2021 205 2051 226
rect 2071 335 2101 355
rect 2071 226 2078 335
rect 2095 226 2101 335
rect 2071 205 2101 226
rect 2121 335 2151 355
rect 2121 226 2128 335
rect 2145 226 2151 335
rect 2219 256 2225 356
rect 2243 256 2249 356
rect 2219 244 2249 256
rect 2309 356 2339 369
rect 2309 256 2315 356
rect 2333 256 2339 356
rect 2309 244 2339 256
rect 2399 356 2429 369
rect 2399 256 2405 356
rect 2423 256 2429 356
rect 2399 244 2429 256
rect 2489 356 2519 369
rect 2489 256 2495 356
rect 2513 256 2519 356
rect 2489 244 2519 256
rect 2579 356 2609 369
rect 2579 256 2585 356
rect 2603 256 2609 356
rect 2579 244 2609 256
rect 2669 356 2699 369
rect 2669 256 2675 356
rect 2693 256 2699 356
rect 2669 244 2699 256
rect 2759 356 2789 369
rect 2759 256 2765 356
rect 2783 256 2789 356
rect 2759 244 2789 256
rect 2849 356 2879 369
rect 2849 256 2855 356
rect 2873 256 2879 356
rect 2849 244 2879 256
rect 2939 356 2969 369
rect 2939 256 2945 356
rect 2963 256 2969 356
rect 2939 244 2969 256
rect 3029 356 3059 369
rect 3029 256 3035 356
rect 3053 256 3059 356
rect 3029 244 3059 256
rect 3119 356 3149 369
rect 3119 256 3125 356
rect 3143 256 3149 356
rect 3119 244 3149 256
rect 3209 356 3239 369
rect 3209 256 3215 356
rect 3233 256 3239 356
rect 3209 244 3239 256
rect 3299 356 3329 369
rect 3299 256 3305 356
rect 3323 256 3329 356
rect 3299 244 3329 256
rect 3389 356 3419 369
rect 3389 256 3395 356
rect 3413 256 3419 356
rect 3389 244 3419 256
rect 3479 356 3509 369
rect 3479 256 3485 356
rect 3503 256 3509 356
rect 3479 244 3509 256
rect 3569 356 3599 369
rect 3569 256 3575 356
rect 3593 256 3599 356
rect 3569 244 3599 256
rect 3659 356 3689 369
rect 3659 256 3665 356
rect 3683 256 3689 356
rect 3659 244 3689 256
rect 3729 356 3759 369
rect 3729 256 3735 356
rect 3753 256 3759 356
rect 3729 244 3759 256
rect 3819 356 3849 369
rect 3819 256 3825 356
rect 3843 256 3849 356
rect 3819 244 3849 256
rect 3909 356 3939 369
rect 3909 256 3915 356
rect 3933 256 3939 356
rect 3909 244 3939 256
rect 3999 356 4029 369
rect 3999 256 4005 356
rect 4023 256 4029 356
rect 3999 244 4029 256
rect 4089 356 4119 369
rect 4089 256 4095 356
rect 4113 256 4119 356
rect 4089 244 4119 256
rect 4179 356 4209 369
rect 4179 256 4185 356
rect 4203 256 4209 356
rect 4179 244 4209 256
rect 4269 356 4299 369
rect 4269 256 4275 356
rect 4293 256 4299 356
rect 4269 244 4299 256
rect 4359 356 4389 369
rect 4359 256 4365 356
rect 4383 256 4389 356
rect 4359 244 4389 256
rect 4449 356 4479 369
rect 4449 256 4455 356
rect 4473 256 4479 356
rect 4449 244 4479 256
rect 4539 356 4569 369
rect 4539 256 4545 356
rect 4563 256 4569 356
rect 4539 244 4569 256
rect 4629 356 4659 369
rect 4629 256 4635 356
rect 4653 256 4659 356
rect 4629 244 4659 256
rect 4719 356 4749 369
rect 4719 256 4725 356
rect 4743 256 4749 356
rect 4719 244 4749 256
rect 4809 356 4839 369
rect 4809 256 4815 356
rect 4833 256 4839 356
rect 4809 244 4839 256
rect 4899 356 4929 369
rect 4899 256 4905 356
rect 4923 256 4929 356
rect 4899 244 4929 256
rect 4989 356 5019 369
rect 4989 256 4995 356
rect 5013 256 5019 356
rect 4989 244 5019 256
rect 5079 356 5109 369
rect 5079 256 5085 356
rect 5103 256 5109 356
rect 5079 244 5109 256
rect 5169 356 5199 369
rect 5169 256 5175 356
rect 5193 256 5199 356
rect 5169 244 5199 256
rect 2121 205 2151 226
<< ndiffc >>
rect -677 463 -660 563
rect -607 463 -590 563
rect -537 463 -520 563
rect -467 463 -450 563
rect -397 463 -380 563
rect -327 463 -310 563
rect -209 478 -191 542
rect -139 478 -121 542
rect -607 130 -589 196
rect -437 130 -419 196
rect -282 92 -265 261
rect -212 92 -195 261
rect -142 92 -125 261
rect 131 58 149 106
rect 221 58 239 106
rect 311 58 329 106
rect 401 58 419 106
rect 491 58 509 106
rect 581 58 599 106
rect 671 58 689 106
rect 761 58 779 106
rect 851 58 869 106
rect 1271 58 1289 106
rect 1361 58 1379 106
rect 1451 58 1469 106
rect 1541 58 1559 106
rect 1631 58 1649 106
rect 1721 58 1739 106
rect 1811 58 1829 106
rect 1901 58 1919 106
rect 1991 58 2009 106
rect 2225 51 2243 151
rect 2315 51 2333 151
rect 2405 51 2423 151
rect 2495 51 2513 151
rect 2585 51 2603 151
rect 2675 51 2693 151
rect 2765 51 2783 151
rect 2855 51 2873 151
rect 2945 51 2963 151
rect 3035 51 3053 151
rect 3125 51 3143 151
rect 3215 51 3233 151
rect 3305 51 3323 151
rect 3395 51 3413 151
rect 3485 51 3503 151
rect 3575 51 3593 151
rect 3665 51 3683 151
rect 3735 51 3753 151
rect 3825 51 3843 151
rect 3915 51 3933 151
rect 4005 51 4023 151
rect 4095 51 4113 151
rect 4185 51 4203 151
rect 4275 51 4293 151
rect 4365 51 4383 151
rect 4455 51 4473 151
rect 4545 51 4563 151
rect 4635 51 4653 151
rect 4725 51 4743 151
rect 4815 51 4833 151
rect 4905 51 4923 151
rect 4995 51 5013 151
rect 5085 51 5103 151
rect 5175 51 5193 151
<< pdiffc >>
rect 40 449 61 582
rect 120 449 141 582
rect 200 449 221 582
rect 280 449 301 582
rect 360 449 381 582
rect 440 449 461 582
rect 520 449 541 582
rect 600 449 621 582
rect 680 449 701 582
rect 760 449 781 582
rect 840 449 861 582
rect 920 449 941 582
rect 1000 449 1021 582
rect 1080 449 1101 582
rect 1160 449 1181 582
rect 1240 449 1261 582
rect 1320 449 1341 582
rect 1400 449 1421 582
rect 1480 449 1501 582
rect 1560 449 1581 582
rect 1640 449 1661 582
rect 1720 449 1741 582
rect 1800 449 1821 582
rect 1880 449 1901 582
rect 1960 449 1981 582
rect 2040 449 2061 582
rect 2120 449 2141 582
rect 2225 471 2243 571
rect 2315 471 2333 571
rect 2405 471 2423 571
rect 2495 471 2513 571
rect 2585 471 2603 571
rect 2675 471 2693 571
rect 2765 471 2783 571
rect 2855 471 2873 571
rect 2945 471 2963 571
rect 3035 471 3053 571
rect 3125 471 3143 571
rect 3215 471 3233 571
rect 3305 471 3323 571
rect 3395 471 3413 571
rect 3485 471 3503 571
rect 3575 471 3593 571
rect 3665 471 3683 571
rect 3735 471 3753 571
rect 3825 471 3843 571
rect 3915 471 3933 571
rect 4005 471 4023 571
rect 4095 471 4113 571
rect 4185 471 4203 571
rect 4275 471 4293 571
rect 4365 471 4383 571
rect 4455 471 4473 571
rect 4545 471 4563 571
rect 4635 471 4653 571
rect 4725 471 4743 571
rect 4815 471 4833 571
rect 4905 471 4923 571
rect 4995 471 5013 571
rect 5085 471 5103 571
rect 5175 471 5193 571
rect 28 226 45 335
rect 78 226 95 335
rect 128 226 145 335
rect 178 226 195 335
rect 228 226 245 335
rect 278 226 295 335
rect 328 226 345 335
rect 378 226 395 335
rect 428 226 445 335
rect 478 226 495 335
rect 528 226 545 335
rect 578 226 595 335
rect 628 226 645 335
rect 678 226 695 335
rect 728 226 745 335
rect 778 226 795 335
rect 828 226 845 335
rect 878 226 895 335
rect 928 226 945 335
rect 978 226 995 335
rect 1028 226 1045 335
rect 1128 226 1145 335
rect 1178 226 1195 335
rect 1228 226 1245 335
rect 1278 226 1295 335
rect 1328 226 1345 335
rect 1378 226 1395 335
rect 1428 226 1445 335
rect 1478 226 1495 335
rect 1528 226 1545 335
rect 1578 226 1595 335
rect 1628 226 1645 335
rect 1678 226 1695 335
rect 1728 226 1745 335
rect 1778 226 1795 335
rect 1828 226 1845 335
rect 1878 226 1895 335
rect 1928 226 1945 335
rect 1978 226 1995 335
rect 2028 226 2045 335
rect 2078 226 2095 335
rect 2128 226 2145 335
rect 2225 256 2243 356
rect 2315 256 2333 356
rect 2405 256 2423 356
rect 2495 256 2513 356
rect 2585 256 2603 356
rect 2675 256 2693 356
rect 2765 256 2783 356
rect 2855 256 2873 356
rect 2945 256 2963 356
rect 3035 256 3053 356
rect 3125 256 3143 356
rect 3215 256 3233 356
rect 3305 256 3323 356
rect 3395 256 3413 356
rect 3485 256 3503 356
rect 3575 256 3593 356
rect 3665 256 3683 356
rect 3735 256 3753 356
rect 3825 256 3843 356
rect 3915 256 3933 356
rect 4005 256 4023 356
rect 4095 256 4113 356
rect 4185 256 4203 356
rect 4275 256 4293 356
rect 4365 256 4383 356
rect 4455 256 4473 356
rect 4545 256 4563 356
rect 4635 256 4653 356
rect 4725 256 4743 356
rect 4815 256 4833 356
rect 4905 256 4923 356
rect 4995 256 5013 356
rect 5085 256 5103 356
rect 5175 256 5193 356
<< psubdiff >>
rect -304 550 -252 579
rect -304 535 -215 550
rect -304 485 -287 535
rect -231 485 -215 535
rect -304 470 -215 485
rect -304 449 -252 470
rect -349 214 -289 276
rect -413 190 -289 214
rect -413 140 -357 190
rect -330 140 -289 190
rect -413 114 -289 140
rect -349 76 -289 114
rect 875 45 914 120
rect 1226 45 1265 120
rect 3689 39 3729 164
<< nsubdiff >>
rect 2150 584 2191 591
rect 2150 459 2219 584
rect 3689 459 3729 584
rect 2150 441 2191 459
rect 1051 205 1121 355
rect 3689 244 3729 369
<< psubdiffcont >>
rect -287 485 -231 535
rect -357 140 -330 190
<< poly >>
rect 70 600 2110 624
rect 3680 609 3728 635
rect -654 579 -614 597
rect -584 579 -544 597
rect -514 579 -474 597
rect -444 579 -404 597
rect -374 579 -334 597
rect 70 591 110 600
rect 150 591 190 600
rect 230 591 270 600
rect 310 591 350 600
rect 390 591 430 600
rect 470 591 510 600
rect 550 591 590 600
rect 630 591 670 600
rect 710 591 750 600
rect 790 591 830 600
rect 870 591 910 600
rect 950 591 990 600
rect 1030 591 1070 600
rect 1110 591 1150 600
rect 1190 591 1230 600
rect 1270 591 1310 600
rect 1350 591 1390 600
rect 1430 591 1470 600
rect 1510 591 1550 600
rect 1590 591 1630 600
rect 1670 591 1710 600
rect 1750 591 1790 600
rect 1830 591 1870 600
rect 1910 591 1950 600
rect 1990 591 2030 600
rect 2070 591 2110 600
rect 2249 594 5170 609
rect -185 550 -145 565
rect -654 429 -614 449
rect -584 429 -544 449
rect -514 429 -474 449
rect -444 429 -404 449
rect -374 429 -334 449
rect -654 398 -334 429
rect -185 443 -145 470
rect -185 426 -174 443
rect -156 426 -145 443
rect 2249 584 2309 594
rect 2339 584 2399 594
rect 2429 584 2489 594
rect 2519 584 2579 594
rect 2609 584 2669 594
rect 2699 584 2759 594
rect 2789 584 2849 594
rect 2879 584 2939 594
rect 2969 584 3029 594
rect 3059 584 3119 594
rect 3149 584 3209 594
rect 3239 584 3299 594
rect 3329 584 3389 594
rect 3419 584 3479 594
rect 3509 584 3569 594
rect 3599 584 3659 594
rect 3759 584 3819 594
rect 3849 584 3909 594
rect 3939 584 3999 594
rect 4029 584 4089 594
rect 4119 584 4179 594
rect 4209 584 4269 594
rect 4299 584 4359 594
rect 4389 584 4449 594
rect 4479 584 4539 594
rect 4569 584 4629 594
rect 4659 584 4719 594
rect 4749 584 4809 594
rect 4839 584 4899 594
rect 4929 584 4989 594
rect 5019 584 5079 594
rect 5109 584 5169 594
rect 2249 445 2309 459
rect 2339 445 2399 459
rect 2429 445 2489 459
rect 2519 445 2579 459
rect 2609 445 2669 459
rect 2699 445 2759 459
rect 2789 445 2849 459
rect 2879 445 2939 459
rect 2969 445 3029 459
rect 3059 445 3119 459
rect 3149 445 3209 459
rect 3239 445 3299 459
rect 3329 445 3389 459
rect 3419 445 3479 459
rect 3509 445 3569 459
rect 3599 445 3659 459
rect 3759 445 3819 459
rect 3849 445 3909 459
rect 3939 445 3999 459
rect 4029 445 4089 459
rect 4119 445 4179 459
rect 4209 445 4269 459
rect 4299 445 4359 459
rect 4389 445 4449 459
rect 4479 445 4539 459
rect 4569 445 4629 459
rect 4659 445 4719 459
rect 4749 445 4809 459
rect 4839 445 4899 459
rect 4929 445 4989 459
rect 5019 445 5079 459
rect 5109 445 5169 459
rect 70 432 110 441
rect -185 418 -145 426
rect -21 416 111 432
rect 150 426 190 441
rect 230 426 270 441
rect 310 426 350 441
rect 390 426 430 441
rect 470 426 510 441
rect 550 426 590 441
rect 630 426 670 441
rect 710 426 750 441
rect 790 426 830 441
rect 870 426 910 441
rect 950 426 990 441
rect 1030 426 1070 441
rect 1110 426 1150 441
rect 1190 426 1230 441
rect 1270 426 1310 441
rect 1350 426 1390 441
rect 1430 426 1470 441
rect 1510 426 1550 441
rect 1590 426 1630 441
rect 1670 426 1710 441
rect 1750 426 1790 441
rect 1830 426 1870 441
rect 1910 426 1950 441
rect 1990 426 2030 441
rect 2070 426 2110 441
rect -654 330 -625 398
rect -670 317 -609 330
rect -670 296 -651 317
rect -627 296 -609 317
rect -670 283 -609 296
rect -419 319 -364 333
rect -419 296 -403 319
rect -379 314 -364 319
rect -379 296 -149 314
rect -419 295 -149 296
rect -419 294 -219 295
rect -419 282 -364 294
rect -259 276 -219 294
rect -189 276 -149 295
rect -553 243 -473 251
rect -553 214 -538 243
rect -485 214 -473 243
rect -553 173 -473 214
rect -553 116 -473 153
rect -21 162 -3 416
rect 51 364 1021 381
rect 51 355 71 364
rect 101 355 121 364
rect 151 355 171 364
rect 201 355 221 364
rect 251 355 271 364
rect 301 355 321 364
rect 351 355 371 364
rect 401 355 421 364
rect 451 355 471 364
rect 501 355 521 364
rect 551 355 571 364
rect 601 355 621 364
rect 651 355 671 364
rect 701 355 721 364
rect 751 355 771 364
rect 801 355 821 364
rect 851 355 871 364
rect 901 355 921 364
rect 951 355 971 364
rect 1001 355 1021 364
rect 1151 363 2121 380
rect 2249 369 2309 383
rect 2339 369 2399 383
rect 2429 369 2489 383
rect 2519 369 2579 383
rect 2609 369 2669 383
rect 2699 369 2759 383
rect 2789 369 2849 383
rect 2879 369 2939 383
rect 2969 369 3029 383
rect 3059 369 3119 383
rect 3149 369 3209 383
rect 3239 369 3299 383
rect 3329 369 3389 383
rect 3419 369 3479 383
rect 3509 369 3569 383
rect 3599 369 3659 383
rect 3759 369 3819 383
rect 3849 369 3909 383
rect 3939 369 3999 383
rect 4029 369 4089 383
rect 4119 369 4179 383
rect 4209 369 4269 383
rect 4299 369 4359 383
rect 4389 369 4449 383
rect 4479 369 4539 383
rect 4569 369 4629 383
rect 4659 369 4719 383
rect 4749 369 4809 383
rect 4839 369 4899 383
rect 4929 369 4989 383
rect 5019 369 5079 383
rect 5109 369 5169 383
rect 1151 355 1171 363
rect 1201 355 1221 363
rect 1251 355 1271 363
rect 1301 355 1321 363
rect 1351 355 1371 363
rect 1401 355 1421 363
rect 1451 355 1471 363
rect 1501 355 1521 363
rect 1551 355 1571 363
rect 1601 355 1621 363
rect 1651 355 1671 363
rect 1701 355 1721 363
rect 1751 355 1771 363
rect 1801 355 1821 363
rect 1851 355 1871 363
rect 1901 355 1921 363
rect 1951 355 1971 363
rect 2001 355 2021 363
rect 2051 355 2071 363
rect 2101 355 2121 363
rect 2249 235 2309 244
rect 2339 235 2399 244
rect 2429 235 2489 244
rect 2519 235 2579 244
rect 2609 235 2669 244
rect 2699 235 2759 244
rect 2789 235 2849 244
rect 2879 235 2939 244
rect 2969 235 3029 244
rect 3059 235 3119 244
rect 3149 235 3209 244
rect 3239 235 3299 244
rect 3329 235 3389 244
rect 3419 235 3479 244
rect 3509 235 3569 244
rect 3599 235 3659 244
rect 3759 235 3819 244
rect 3849 235 3909 244
rect 3939 235 3999 244
rect 4029 235 4089 244
rect 4119 235 4179 244
rect 4209 235 4269 244
rect 4299 235 4359 244
rect 4389 235 4449 244
rect 4479 235 4539 244
rect 4569 235 4629 244
rect 4659 235 4719 244
rect 4749 235 4809 244
rect 4839 235 4899 244
rect 4929 235 4989 244
rect 5019 235 5079 244
rect 5109 235 5169 244
rect 2249 220 5170 235
rect 3687 215 3733 220
rect 51 192 71 205
rect 101 192 121 205
rect 151 192 171 205
rect 201 192 221 205
rect 251 192 271 205
rect 301 192 321 205
rect 351 192 371 205
rect 401 192 421 205
rect 451 192 471 205
rect 501 192 521 205
rect 551 192 571 205
rect 601 192 621 205
rect 651 192 671 205
rect 701 192 721 205
rect 751 192 771 205
rect 801 192 821 205
rect 851 192 871 205
rect 901 192 921 205
rect 951 192 971 205
rect -21 153 17 162
rect -21 134 -12 153
rect 7 134 17 153
rect -21 126 17 134
rect 1001 133 1021 205
rect 1151 133 1171 205
rect 1201 192 1221 205
rect 1251 192 1271 205
rect 1301 192 1321 205
rect 1351 192 1371 205
rect 1401 192 1421 205
rect 1451 192 1471 205
rect 1501 192 1521 205
rect 1551 192 1571 205
rect 1601 192 1621 205
rect 1651 192 1671 205
rect 1701 192 1721 205
rect 1751 192 1771 205
rect 1801 192 1821 205
rect 1851 192 1871 205
rect 1901 192 1921 205
rect 1951 192 1971 205
rect 2001 192 2021 205
rect 2051 192 2071 205
rect 2101 192 2121 205
rect 3687 192 3699 215
rect 3721 192 3733 215
rect 3687 182 3733 192
rect 2249 164 2309 178
rect 2339 164 2399 178
rect 2429 164 2489 178
rect 2519 164 2579 178
rect 2609 164 2669 178
rect 2699 164 2759 178
rect 2789 164 2849 178
rect 2879 164 2939 178
rect 2969 164 3029 178
rect 3059 164 3119 178
rect 3149 164 3209 178
rect 3239 164 3299 178
rect 3329 164 3389 178
rect 3419 164 3479 178
rect 3509 164 3569 178
rect 3599 164 3659 178
rect 3759 164 3819 178
rect 3849 164 3909 178
rect 3939 164 3999 178
rect 4029 164 4089 178
rect 4119 164 4179 178
rect 4209 164 4269 178
rect 4299 164 4359 178
rect 4389 164 4449 178
rect 4479 164 4539 178
rect 4569 164 4629 178
rect 4659 164 4719 178
rect 4749 164 4809 178
rect 4839 164 4899 178
rect 4929 164 4989 178
rect 5019 164 5079 178
rect 5109 164 5169 178
rect 155 120 215 133
rect 245 120 305 133
rect 335 120 395 133
rect 425 120 485 133
rect 515 120 575 133
rect 605 120 665 133
rect 695 120 755 133
rect 785 120 845 133
rect 993 125 1031 133
rect -259 53 -219 76
rect -189 53 -149 76
rect 42 46 78 55
rect 42 28 51 46
rect 69 37 78 46
rect 993 108 1002 125
rect 1022 108 1031 125
rect 993 101 1031 108
rect 1143 125 1181 133
rect 1143 108 1152 125
rect 1172 108 1181 125
rect 1295 120 1355 133
rect 1385 120 1445 133
rect 1475 120 1535 133
rect 1565 120 1625 133
rect 1655 120 1715 133
rect 1745 120 1805 133
rect 1835 120 1895 133
rect 1925 120 1985 133
rect 1143 101 1181 108
rect 155 37 215 45
rect 245 37 305 45
rect 335 37 395 45
rect 425 37 485 45
rect 515 37 575 45
rect 605 37 665 45
rect 695 37 755 45
rect 785 37 845 45
rect 1295 37 1355 45
rect 1385 37 1445 45
rect 1475 37 1535 45
rect 1565 37 1625 45
rect 1655 37 1715 45
rect 1745 37 1805 45
rect 1835 37 1895 45
rect 1925 37 1985 45
rect 5224 41 5257 49
rect 69 28 1985 37
rect 2249 29 2309 39
rect 2339 29 2399 39
rect 2429 29 2489 39
rect 2519 29 2579 39
rect 2609 29 2669 39
rect 2699 29 2759 39
rect 2789 29 2849 39
rect 2879 29 2939 39
rect 2969 29 3029 39
rect 3059 29 3119 39
rect 3149 29 3209 39
rect 3239 29 3299 39
rect 3329 29 3389 39
rect 3419 29 3479 39
rect 3509 29 3569 39
rect 3599 29 3659 39
rect 3759 29 3819 39
rect 3849 29 3909 39
rect 3939 29 3999 39
rect 4029 29 4089 39
rect 4119 29 4179 39
rect 4209 29 4269 39
rect 4299 29 4359 39
rect 4389 29 4449 39
rect 4479 29 4539 39
rect 4569 29 4629 39
rect 4659 29 4719 39
rect 4749 29 4809 39
rect 4839 29 4899 39
rect 4929 29 4989 39
rect 5019 29 5079 39
rect 5109 29 5169 39
rect 5224 29 5232 41
rect 42 22 1985 28
rect 2248 23 5232 29
rect 5250 23 5257 41
rect 42 20 78 22
rect 2248 14 5257 23
<< polycont >>
rect -174 426 -156 443
rect -651 296 -627 317
rect -403 296 -379 319
rect -538 214 -485 243
rect -12 134 7 153
rect 3699 192 3721 215
rect 51 28 69 46
rect 1002 108 1022 125
rect 1152 108 1172 125
rect 5232 23 5250 41
<< locali >>
rect -508 643 -444 653
rect -508 620 -489 643
rect -464 620 -444 643
rect 1213 642 1284 653
rect 1213 632 1236 642
rect 113 620 1236 632
rect 1262 632 1284 642
rect 2826 644 2899 653
rect 1262 620 2067 632
rect 2826 624 2849 644
rect -613 601 -305 620
rect -683 563 -655 579
rect -683 463 -677 563
rect -660 463 -655 563
rect -683 420 -655 463
rect -613 563 -585 601
rect -613 463 -607 563
rect -590 463 -585 563
rect -613 449 -585 463
rect -543 563 -515 579
rect -543 463 -537 563
rect -520 463 -515 563
rect -543 420 -515 463
rect -473 563 -445 601
rect -333 579 -305 601
rect 113 610 2067 620
rect 33 582 67 591
rect -473 463 -467 563
rect -450 463 -445 563
rect -473 449 -445 463
rect -403 563 -375 579
rect -403 463 -397 563
rect -380 463 -375 563
rect -403 420 -375 463
rect -333 563 -252 579
rect -333 463 -327 563
rect -310 550 -252 563
rect -310 542 -186 550
rect -310 535 -209 542
rect -310 485 -287 535
rect -231 485 -209 535
rect -310 478 -209 485
rect -191 478 -186 542
rect -310 470 -186 478
rect -144 542 -116 550
rect -144 478 -139 542
rect -121 478 -116 542
rect -310 463 -252 470
rect -333 449 -252 463
rect -144 453 -116 478
rect -684 400 -375 420
rect -218 443 -116 453
rect -218 426 -174 443
rect -156 426 -116 443
rect -218 418 -116 426
rect 33 449 40 582
rect 61 449 67 582
rect -542 348 -515 400
rect -218 381 -189 418
rect 33 408 67 449
rect 113 582 147 610
rect 113 449 120 582
rect 141 449 147 582
rect 113 441 147 449
rect 193 582 227 591
rect 193 449 200 582
rect 221 449 227 582
rect 193 408 227 449
rect 273 582 307 610
rect 273 449 280 582
rect 301 449 307 582
rect 273 441 307 449
rect 353 582 387 591
rect 353 449 360 582
rect 381 449 387 582
rect 353 408 387 449
rect 433 582 467 610
rect 433 449 440 582
rect 461 449 467 582
rect 433 441 467 449
rect 513 582 547 591
rect 513 449 520 582
rect 541 449 547 582
rect 513 408 547 449
rect 593 582 627 610
rect 593 449 600 582
rect 621 449 627 582
rect 593 441 627 449
rect 673 582 707 591
rect 673 449 680 582
rect 701 449 707 582
rect 673 408 707 449
rect 753 582 787 610
rect 753 449 760 582
rect 781 449 787 582
rect 753 441 787 449
rect 833 582 867 591
rect 833 449 840 582
rect 861 449 867 582
rect 833 408 867 449
rect 913 582 947 610
rect 913 449 920 582
rect 941 449 947 582
rect 913 441 947 449
rect 993 582 1027 591
rect 993 449 1000 582
rect 1021 449 1027 582
rect 993 408 1027 449
rect 1073 582 1107 610
rect 1073 449 1080 582
rect 1101 449 1107 582
rect 1073 441 1107 449
rect 1153 582 1187 591
rect 1153 449 1160 582
rect 1181 449 1187 582
rect 1153 408 1187 449
rect 1233 582 1267 610
rect 1233 449 1240 582
rect 1261 449 1267 582
rect 1233 441 1267 449
rect 1313 582 1347 591
rect 1313 449 1320 582
rect 1341 449 1347 582
rect 1313 408 1347 449
rect 1393 582 1427 610
rect 1393 449 1400 582
rect 1421 449 1427 582
rect 1393 441 1427 449
rect 1473 582 1507 591
rect 1473 449 1480 582
rect 1501 449 1507 582
rect 1473 408 1507 449
rect 1553 582 1587 610
rect 1553 449 1560 582
rect 1581 449 1587 582
rect 1553 441 1587 449
rect 1633 582 1667 591
rect 1633 449 1640 582
rect 1661 449 1667 582
rect 1633 408 1667 449
rect 1713 582 1747 610
rect 1713 449 1720 582
rect 1741 449 1747 582
rect 1713 441 1747 449
rect 1793 582 1827 591
rect 1793 449 1800 582
rect 1821 449 1827 582
rect 1793 408 1827 449
rect 1873 582 1907 610
rect 1873 449 1880 582
rect 1901 449 1907 582
rect 1873 441 1907 449
rect 1953 582 1987 591
rect 1953 449 1960 582
rect 1981 449 1987 582
rect 1953 408 1987 449
rect 2033 582 2067 610
rect 2311 618 2849 624
rect 2876 624 2899 644
rect 4348 644 4400 653
rect 3680 630 3728 635
rect 4348 631 4361 644
rect 2876 618 3597 624
rect 2311 607 3597 618
rect 3680 613 3695 630
rect 3712 613 3728 630
rect 3680 609 3728 613
rect 3821 621 4361 631
rect 4387 631 4400 644
rect 4387 621 5107 631
rect 3821 611 5107 621
rect 2033 449 2040 582
rect 2061 449 2067 582
rect 2033 441 2067 449
rect 2113 582 2147 591
rect 2113 449 2120 582
rect 2141 449 2147 582
rect 2113 408 2147 449
rect 2221 571 2247 584
rect 2221 471 2225 571
rect 2243 471 2247 571
rect 2221 429 2247 471
rect 2311 571 2337 607
rect 2311 471 2315 571
rect 2333 471 2337 571
rect 2311 459 2337 471
rect 2401 571 2427 584
rect 2401 471 2405 571
rect 2423 471 2427 571
rect 2401 429 2427 471
rect 2491 571 2517 607
rect 2491 471 2495 571
rect 2513 471 2517 571
rect 2491 459 2517 471
rect 2581 571 2607 584
rect 2581 471 2585 571
rect 2603 471 2607 571
rect 2581 429 2607 471
rect 2671 571 2697 607
rect 2671 471 2675 571
rect 2693 471 2697 571
rect 2671 459 2697 471
rect 2761 571 2787 584
rect 2761 471 2765 571
rect 2783 471 2787 571
rect 2761 429 2787 471
rect 2851 571 2877 607
rect 2851 471 2855 571
rect 2873 471 2877 571
rect 2851 459 2877 471
rect 2941 571 2967 584
rect 2941 471 2945 571
rect 2963 471 2967 571
rect 2941 429 2967 471
rect 3031 571 3057 607
rect 3031 471 3035 571
rect 3053 471 3057 571
rect 3031 459 3057 471
rect 3121 571 3147 584
rect 3121 471 3125 571
rect 3143 471 3147 571
rect 3121 429 3147 471
rect 3211 571 3237 607
rect 3211 471 3215 571
rect 3233 471 3237 571
rect 3211 459 3237 471
rect 3301 571 3327 584
rect 3301 471 3305 571
rect 3323 471 3327 571
rect 3301 429 3327 471
rect 3391 571 3417 607
rect 3391 471 3395 571
rect 3413 471 3417 571
rect 3391 459 3417 471
rect 3481 571 3507 584
rect 3481 471 3485 571
rect 3503 471 3507 571
rect 3481 429 3507 471
rect 3571 571 3597 607
rect 3571 471 3575 571
rect 3593 471 3597 571
rect 3571 459 3597 471
rect 3661 571 3687 584
rect 3661 471 3665 571
rect 3683 471 3687 571
rect 3661 429 3687 471
rect 23 385 2149 408
rect -218 363 -139 381
rect -542 332 -480 348
rect -218 334 -183 363
rect -153 334 -139 363
rect -670 317 -609 330
rect -670 296 -651 317
rect -627 296 -609 317
rect -670 283 -609 296
rect -542 308 -522 332
rect -497 308 -480 332
rect -542 296 -480 308
rect -419 319 -364 333
rect -419 296 -403 319
rect -379 296 -364 319
rect -542 251 -515 296
rect -419 282 -364 296
rect -218 323 -139 334
rect 23 335 49 385
rect -288 261 -260 276
rect -613 243 -470 251
rect -613 230 -538 243
rect -612 196 -584 230
rect -553 214 -538 230
rect -485 214 -470 243
rect -553 206 -470 214
rect -612 130 -607 196
rect -589 130 -584 196
rect -612 114 -584 130
rect -442 196 -414 214
rect -442 130 -437 196
rect -419 180 -414 196
rect -368 190 -321 201
rect -368 180 -357 190
rect -419 145 -357 180
rect -419 130 -414 145
rect -442 114 -414 130
rect -368 140 -357 145
rect -330 180 -321 190
rect -288 180 -282 261
rect -330 145 -282 180
rect -330 140 -321 145
rect -368 129 -321 140
rect -288 92 -282 145
rect -265 92 -260 261
rect -288 54 -260 92
rect -218 274 -189 323
rect -218 261 -190 274
rect -218 92 -212 261
rect -195 92 -190 261
rect -218 76 -190 92
rect -148 261 -120 276
rect -148 92 -142 261
rect -125 92 -120 261
rect 23 226 28 335
rect 45 226 49 335
rect 23 205 49 226
rect 73 335 99 355
rect 73 226 78 335
rect 95 226 99 335
rect 73 173 99 226
rect 123 335 149 385
rect 123 226 128 335
rect 145 226 149 335
rect 123 205 149 226
rect 173 335 199 355
rect 173 226 178 335
rect 195 226 199 335
rect 173 173 199 226
rect 223 335 249 385
rect 223 226 228 335
rect 245 226 249 335
rect 223 205 249 226
rect 273 335 299 355
rect 273 226 278 335
rect 295 226 299 335
rect 273 173 299 226
rect 323 335 349 385
rect 323 226 328 335
rect 345 226 349 335
rect 323 205 349 226
rect 373 335 399 355
rect 373 226 378 335
rect 395 226 399 335
rect 373 173 399 226
rect 423 335 449 385
rect 423 226 428 335
rect 445 226 449 335
rect 423 205 449 226
rect 473 335 499 355
rect 473 226 478 335
rect 495 226 499 335
rect 473 173 499 226
rect 523 335 549 385
rect 523 226 528 335
rect 545 226 549 335
rect 523 205 549 226
rect 573 335 599 355
rect 573 226 578 335
rect 595 226 599 335
rect 573 173 599 226
rect 623 335 649 385
rect 623 226 628 335
rect 645 226 649 335
rect 623 205 649 226
rect 673 335 699 355
rect 673 226 678 335
rect 695 226 699 335
rect 673 173 699 226
rect 723 335 749 385
rect 723 226 728 335
rect 745 226 749 335
rect 723 205 749 226
rect 773 335 799 355
rect 773 226 778 335
rect 795 226 799 335
rect 773 173 799 226
rect 823 335 849 385
rect 823 226 828 335
rect 845 226 849 335
rect 823 205 849 226
rect 873 335 899 355
rect 873 226 878 335
rect 895 226 899 335
rect 873 173 899 226
rect 923 335 949 385
rect 923 226 928 335
rect 945 226 949 335
rect 923 205 949 226
rect 973 335 999 355
rect 973 226 978 335
rect 995 226 999 335
rect 973 173 999 226
rect 1023 335 1049 385
rect 1023 226 1028 335
rect 1045 226 1049 335
rect 1023 205 1049 226
rect 1123 335 1149 385
rect 1123 226 1128 335
rect 1145 226 1149 335
rect 1123 209 1149 226
rect 1173 335 1199 355
rect 1173 226 1178 335
rect 1195 226 1199 335
rect -21 153 17 162
rect -21 134 -12 153
rect 7 134 17 153
rect 73 150 999 173
rect 1173 175 1199 226
rect 1223 335 1249 385
rect 1223 226 1228 335
rect 1245 226 1249 335
rect 1223 205 1249 226
rect 1273 335 1299 355
rect 1273 226 1278 335
rect 1295 226 1299 335
rect 1273 175 1299 226
rect 1323 335 1349 385
rect 1323 226 1328 335
rect 1345 226 1349 335
rect 1323 205 1349 226
rect 1373 335 1399 355
rect 1373 226 1378 335
rect 1395 226 1399 335
rect 1373 175 1399 226
rect 1423 335 1449 385
rect 1423 226 1428 335
rect 1445 226 1449 335
rect 1423 205 1449 226
rect 1473 335 1499 355
rect 1473 226 1478 335
rect 1495 226 1499 335
rect 1473 175 1499 226
rect 1523 335 1549 385
rect 1523 226 1528 335
rect 1545 226 1549 335
rect 1523 205 1549 226
rect 1573 335 1599 355
rect 1573 226 1578 335
rect 1595 226 1599 335
rect 1573 175 1599 226
rect 1623 335 1649 385
rect 1623 226 1628 335
rect 1645 226 1649 335
rect 1623 205 1649 226
rect 1673 335 1699 355
rect 1673 226 1678 335
rect 1695 226 1699 335
rect 1673 175 1699 226
rect 1723 335 1749 385
rect 1723 226 1728 335
rect 1745 226 1749 335
rect 1723 205 1749 226
rect 1773 335 1799 355
rect 1773 226 1778 335
rect 1795 226 1799 335
rect 1773 175 1799 226
rect 1823 335 1849 385
rect 1823 226 1828 335
rect 1845 226 1849 335
rect 1823 205 1849 226
rect 1873 335 1899 355
rect 1873 226 1878 335
rect 1895 226 1899 335
rect 1873 175 1899 226
rect 1923 335 1949 385
rect 1923 226 1928 335
rect 1945 226 1949 335
rect 1923 205 1949 226
rect 1973 335 1999 355
rect 1973 226 1978 335
rect 1995 226 1999 335
rect 1973 175 1999 226
rect 2023 335 2049 385
rect 2023 226 2028 335
rect 2045 226 2049 335
rect 2023 205 2049 226
rect 2073 335 2099 355
rect 2073 226 2078 335
rect 2095 226 2099 335
rect 2073 175 2099 226
rect 2123 335 2149 385
rect 2123 226 2128 335
rect 2145 226 2149 335
rect 2221 398 3687 429
rect 2221 356 2247 398
rect 2221 256 2225 356
rect 2243 256 2247 356
rect 2221 244 2247 256
rect 2311 356 2337 369
rect 2311 256 2315 356
rect 2333 256 2337 356
rect 2123 205 2149 226
rect 2311 217 2337 256
rect 2401 356 2427 398
rect 2401 256 2405 356
rect 2423 256 2427 356
rect 2401 244 2427 256
rect 2491 356 2517 369
rect 2491 256 2495 356
rect 2513 256 2517 356
rect 2491 217 2517 256
rect 2581 356 2607 398
rect 2581 256 2585 356
rect 2603 256 2607 356
rect 2581 244 2607 256
rect 2671 356 2697 369
rect 2671 256 2675 356
rect 2693 256 2697 356
rect 2671 217 2697 256
rect 2761 356 2787 398
rect 2761 256 2765 356
rect 2783 256 2787 356
rect 2761 244 2787 256
rect 2851 356 2877 369
rect 2851 256 2855 356
rect 2873 256 2877 356
rect 2851 217 2877 256
rect 2941 356 2967 398
rect 2941 256 2945 356
rect 2963 256 2967 356
rect 2941 244 2967 256
rect 3031 356 3057 369
rect 3031 256 3035 356
rect 3053 256 3057 356
rect 3031 217 3057 256
rect 3121 356 3147 398
rect 3121 256 3125 356
rect 3143 256 3147 356
rect 3121 244 3147 256
rect 3211 356 3237 369
rect 3211 256 3215 356
rect 3233 256 3237 356
rect 3211 217 3237 256
rect 3301 356 3327 398
rect 3301 256 3305 356
rect 3323 256 3327 356
rect 3301 244 3327 256
rect 3391 356 3417 369
rect 3391 256 3395 356
rect 3413 256 3417 356
rect 3391 217 3417 256
rect 3481 356 3507 398
rect 3481 256 3485 356
rect 3503 256 3507 356
rect 3481 244 3507 256
rect 3571 356 3597 369
rect 3571 256 3575 356
rect 3593 256 3597 356
rect 3571 217 3597 256
rect 3661 356 3687 398
rect 3661 256 3665 356
rect 3683 256 3687 356
rect 3661 244 3687 256
rect 3731 571 3757 584
rect 3731 471 3735 571
rect 3753 471 3757 571
rect 3731 430 3757 471
rect 3821 571 3847 611
rect 3821 471 3825 571
rect 3843 471 3847 571
rect 3821 459 3847 471
rect 3911 571 3937 584
rect 3911 471 3915 571
rect 3933 471 3937 571
rect 3911 430 3937 471
rect 4001 571 4027 611
rect 4001 471 4005 571
rect 4023 471 4027 571
rect 4001 459 4027 471
rect 4091 571 4117 584
rect 4091 471 4095 571
rect 4113 471 4117 571
rect 4091 430 4117 471
rect 4181 571 4207 611
rect 4181 471 4185 571
rect 4203 471 4207 571
rect 4181 459 4207 471
rect 4271 571 4297 584
rect 4271 471 4275 571
rect 4293 471 4297 571
rect 4271 430 4297 471
rect 4361 571 4387 611
rect 4361 471 4365 571
rect 4383 471 4387 571
rect 4361 459 4387 471
rect 4451 571 4477 584
rect 4451 471 4455 571
rect 4473 471 4477 571
rect 4451 430 4477 471
rect 4541 571 4567 611
rect 4541 471 4545 571
rect 4563 471 4567 571
rect 4541 459 4567 471
rect 4631 571 4657 584
rect 4631 471 4635 571
rect 4653 471 4657 571
rect 4631 430 4657 471
rect 4721 571 4747 611
rect 4721 471 4725 571
rect 4743 471 4747 571
rect 4721 459 4747 471
rect 4811 571 4837 584
rect 4811 471 4815 571
rect 4833 471 4837 571
rect 4811 430 4837 471
rect 4901 571 4927 611
rect 4901 471 4905 571
rect 4923 471 4927 571
rect 4901 459 4927 471
rect 4991 571 5017 584
rect 4991 471 4995 571
rect 5013 471 5017 571
rect 4991 430 5017 471
rect 5081 571 5107 611
rect 5081 471 5085 571
rect 5103 471 5107 571
rect 5081 459 5107 471
rect 5171 571 5197 584
rect 5171 471 5175 571
rect 5193 471 5197 571
rect 5171 430 5197 471
rect 3731 400 5197 430
rect 3731 356 3757 400
rect 3731 256 3735 356
rect 3753 256 3757 356
rect 3731 244 3757 256
rect 3821 356 3847 369
rect 3821 256 3825 356
rect 3843 256 3847 356
rect 1173 150 2099 175
rect 2311 191 3597 217
rect 2221 151 2247 164
rect -21 126 17 134
rect -148 54 -120 92
rect 127 106 153 150
rect 127 58 131 106
rect 149 58 153 106
rect -288 35 -120 54
rect 42 46 78 55
rect -227 26 -176 35
rect -227 2 -213 26
rect -188 2 -176 26
rect 42 28 51 46
rect 69 28 78 46
rect 127 45 153 58
rect 217 106 243 120
rect 217 58 221 106
rect 239 58 243 106
rect 42 20 78 28
rect 217 25 243 58
rect 307 106 333 150
rect 307 58 311 106
rect 329 58 333 106
rect 307 45 333 58
rect 397 106 423 120
rect 397 58 401 106
rect 419 58 423 106
rect 397 25 423 58
rect 487 106 513 150
rect 487 58 491 106
rect 509 58 513 106
rect 487 45 513 58
rect 577 106 603 120
rect 577 58 581 106
rect 599 58 603 106
rect 577 25 603 58
rect 667 106 693 150
rect 667 58 671 106
rect 689 58 693 106
rect 667 45 693 58
rect 757 106 783 120
rect 757 58 761 106
rect 779 58 783 106
rect 757 25 783 58
rect 847 106 873 150
rect 847 96 851 106
rect 847 78 850 96
rect 847 58 851 78
rect 869 58 873 106
rect 993 125 1031 133
rect 993 108 1002 125
rect 1022 108 1031 125
rect 993 101 1031 108
rect 1143 125 1181 133
rect 1143 108 1152 125
rect 1172 108 1181 125
rect 1143 101 1181 108
rect 1267 106 1293 150
rect 847 45 873 58
rect 1267 58 1271 106
rect 1289 58 1293 106
rect 1267 45 1293 58
rect 1357 106 1383 120
rect 1357 58 1361 106
rect 1379 58 1383 106
rect 1357 25 1383 58
rect 1447 106 1473 150
rect 1447 58 1451 106
rect 1469 58 1473 106
rect 1447 45 1473 58
rect 1537 106 1563 120
rect 1537 58 1541 106
rect 1559 58 1563 106
rect 1537 25 1563 58
rect 1627 106 1653 150
rect 1627 58 1631 106
rect 1649 58 1653 106
rect 1627 45 1653 58
rect 1717 106 1743 120
rect 1717 58 1721 106
rect 1739 58 1743 106
rect 1717 25 1743 58
rect 1807 106 1833 150
rect 1807 58 1811 106
rect 1829 58 1833 106
rect 1807 45 1833 58
rect 1897 106 1923 120
rect 1897 58 1901 106
rect 1919 58 1923 106
rect 1897 25 1923 58
rect 1987 106 2013 150
rect 1987 58 1991 106
rect 2009 58 2013 106
rect 1987 45 2013 58
rect 2221 51 2225 151
rect 2243 51 2247 151
rect 217 19 1923 25
rect 217 3 578 19
rect -227 -7 -176 2
rect 553 1 578 3
rect 598 3 1923 19
rect 2221 22 2247 51
rect 2311 151 2337 191
rect 2311 51 2315 151
rect 2333 51 2337 151
rect 2311 39 2337 51
rect 2401 151 2427 164
rect 2401 51 2405 151
rect 2423 51 2427 151
rect 2401 22 2427 51
rect 2491 151 2517 191
rect 2491 51 2495 151
rect 2513 51 2517 151
rect 2491 39 2517 51
rect 2581 151 2607 164
rect 2581 51 2585 151
rect 2603 51 2607 151
rect 2221 21 2427 22
rect 2581 21 2607 51
rect 2671 151 2697 191
rect 2671 51 2675 151
rect 2693 51 2697 151
rect 2671 39 2697 51
rect 2761 151 2787 164
rect 2761 51 2765 151
rect 2783 51 2787 151
rect 2761 21 2787 51
rect 2851 151 2877 191
rect 2851 51 2855 151
rect 2873 51 2877 151
rect 2851 39 2877 51
rect 2941 151 2967 164
rect 2941 51 2945 151
rect 2963 51 2967 151
rect 2941 21 2967 51
rect 3031 151 3057 191
rect 3031 51 3035 151
rect 3053 51 3057 151
rect 3031 39 3057 51
rect 3121 151 3147 164
rect 3121 51 3125 151
rect 3143 51 3147 151
rect 3121 21 3147 51
rect 3211 151 3237 191
rect 3211 51 3215 151
rect 3233 51 3237 151
rect 3211 39 3237 51
rect 3301 151 3327 164
rect 3301 51 3305 151
rect 3323 51 3327 151
rect 3301 21 3327 51
rect 3391 151 3417 191
rect 3391 51 3395 151
rect 3413 51 3417 151
rect 3391 39 3417 51
rect 3481 151 3507 164
rect 3481 51 3485 151
rect 3503 51 3507 151
rect 3481 21 3507 51
rect 3571 151 3597 191
rect 3687 215 3733 227
rect 3687 192 3699 215
rect 3721 192 3733 215
rect 3687 182 3733 192
rect 3821 216 3847 256
rect 3911 356 3937 400
rect 3911 256 3915 356
rect 3933 256 3937 356
rect 3911 244 3937 256
rect 4001 356 4027 369
rect 4001 256 4005 356
rect 4023 256 4027 356
rect 4001 216 4027 256
rect 4091 356 4117 400
rect 4091 256 4095 356
rect 4113 256 4117 356
rect 4091 244 4117 256
rect 4181 356 4207 369
rect 4181 256 4185 356
rect 4203 256 4207 356
rect 4181 216 4207 256
rect 4271 356 4297 400
rect 4271 256 4275 356
rect 4293 256 4297 356
rect 4271 244 4297 256
rect 4361 356 4387 369
rect 4361 256 4365 356
rect 4383 256 4387 356
rect 4361 216 4387 256
rect 4451 356 4477 400
rect 4451 256 4455 356
rect 4473 256 4477 356
rect 4451 244 4477 256
rect 4541 356 4567 369
rect 4541 256 4545 356
rect 4563 256 4567 356
rect 4541 216 4567 256
rect 4631 356 4657 400
rect 4631 256 4635 356
rect 4653 256 4657 356
rect 4631 244 4657 256
rect 4721 356 4747 369
rect 4721 256 4725 356
rect 4743 256 4747 356
rect 4721 216 4747 256
rect 4811 356 4837 400
rect 4811 256 4815 356
rect 4833 256 4837 356
rect 4811 244 4837 256
rect 4901 356 4927 369
rect 4901 256 4905 356
rect 4923 256 4927 356
rect 4901 216 4927 256
rect 4991 356 5017 400
rect 4991 256 4995 356
rect 5013 256 5017 356
rect 4991 244 5017 256
rect 5081 356 5107 369
rect 5081 256 5085 356
rect 5103 256 5107 356
rect 5081 216 5107 256
rect 5171 356 5197 400
rect 5171 256 5175 356
rect 5193 256 5197 356
rect 5171 244 5197 256
rect 3821 190 5107 216
rect 3571 51 3575 151
rect 3593 51 3597 151
rect 3571 39 3597 51
rect 3661 151 3687 164
rect 3661 51 3665 151
rect 3683 51 3687 151
rect 3661 21 3687 51
rect 2221 4 3687 21
rect 3731 151 3757 164
rect 3731 51 3735 151
rect 3753 51 3757 151
rect 3731 21 3757 51
rect 3821 151 3847 190
rect 3821 51 3825 151
rect 3843 51 3847 151
rect 3821 39 3847 51
rect 3911 151 3937 164
rect 3911 51 3915 151
rect 3933 51 3937 151
rect 3911 21 3937 51
rect 4001 151 4027 190
rect 4001 51 4005 151
rect 4023 51 4027 151
rect 4001 39 4027 51
rect 4091 151 4117 164
rect 4091 51 4095 151
rect 4113 51 4117 151
rect 4091 21 4117 51
rect 4181 151 4207 190
rect 4181 51 4185 151
rect 4203 51 4207 151
rect 4181 39 4207 51
rect 4271 151 4297 164
rect 4271 51 4275 151
rect 4293 51 4297 151
rect 4271 21 4297 51
rect 4361 151 4387 190
rect 4361 51 4365 151
rect 4383 51 4387 151
rect 4361 39 4387 51
rect 4451 151 4477 164
rect 4451 51 4455 151
rect 4473 51 4477 151
rect 4451 21 4477 51
rect 4541 151 4567 190
rect 4541 51 4545 151
rect 4563 51 4567 151
rect 4541 39 4567 51
rect 4631 151 4657 164
rect 4631 51 4635 151
rect 4653 51 4657 151
rect 4631 21 4657 51
rect 4721 151 4747 190
rect 4721 51 4725 151
rect 4743 51 4747 151
rect 4721 39 4747 51
rect 4811 151 4837 164
rect 4811 51 4815 151
rect 4833 51 4837 151
rect 4811 21 4837 51
rect 4901 151 4927 190
rect 4901 51 4905 151
rect 4923 51 4927 151
rect 4901 39 4927 51
rect 4991 151 5017 164
rect 4991 51 4995 151
rect 5013 51 5017 151
rect 4991 21 5017 51
rect 5081 151 5107 190
rect 5081 51 5085 151
rect 5103 51 5107 151
rect 5081 39 5107 51
rect 5171 151 5197 164
rect 5171 51 5175 151
rect 5193 51 5197 151
rect 5171 21 5197 51
rect 3731 3 5197 21
rect 5224 41 5257 49
rect 5224 23 5232 41
rect 5250 23 5257 41
rect 5224 14 5257 23
rect 598 1 622 3
rect 553 -6 622 1
<< viali >>
rect -489 620 -464 643
rect 1236 620 1262 642
rect 2849 618 2876 644
rect 3695 613 3712 630
rect 4361 621 4387 644
rect -183 334 -153 363
rect -651 296 -627 317
rect -522 308 -497 332
rect -403 296 -379 319
rect -12 134 7 153
rect 3575 330 3593 348
rect 3575 293 3593 311
rect -213 2 -188 26
rect 51 28 69 46
rect 850 78 851 96
rect 851 78 868 96
rect 1002 108 1022 125
rect 1152 108 1172 125
rect 1991 86 2009 104
rect 2225 83 2243 100
rect 578 1 598 19
rect 3699 192 3721 215
rect 5085 262 5103 281
rect 3735 103 3753 121
rect 3735 66 3753 84
rect 5232 23 5250 41
<< metal1 >>
rect -508 646 -444 653
rect -508 615 -499 646
rect -450 615 -444 646
rect -508 609 -444 615
rect 1206 647 1294 653
rect 1206 609 1218 647
rect 1282 609 1294 647
rect 1206 603 1294 609
rect 2826 645 2899 653
rect 2826 613 2834 645
rect 2891 613 2899 645
rect 4348 649 4400 653
rect 3680 631 3728 635
rect 2826 607 2899 613
rect 3618 630 3728 631
rect 3618 616 3695 630
rect 1151 467 1203 473
rect 1151 431 1157 467
rect 1197 431 1203 467
rect 1151 425 1203 431
rect -197 363 -139 381
rect -541 332 -480 348
rect -197 334 -183 363
rect -153 334 -139 363
rect -670 323 -609 330
rect -670 289 -660 323
rect -618 289 -609 323
rect -541 308 -522 332
rect -497 308 -480 332
rect -541 296 -480 308
rect -419 327 -364 333
rect -670 283 -609 289
rect -523 121 -498 296
rect -419 288 -409 327
rect -372 288 -364 327
rect -197 323 -139 334
rect -419 282 -364 288
rect -188 169 -155 323
rect 1151 192 1172 425
rect 3618 383 3643 616
rect 3680 613 3695 616
rect 3712 613 3728 630
rect 3680 609 3728 613
rect 4348 617 4354 649
rect 4395 617 4400 649
rect 4348 611 4400 617
rect 3571 361 3643 383
rect 3571 348 3597 361
rect 3571 330 3575 348
rect 3593 330 3597 348
rect 3571 311 3597 330
rect 3571 293 3575 311
rect 3593 293 3597 311
rect 3571 279 3597 293
rect 5074 281 5114 296
rect 5074 262 5085 281
rect 5103 280 5114 281
rect 5103 262 5271 280
rect 5074 255 5271 262
rect 5074 249 5114 255
rect 3687 219 3733 227
rect 993 180 1031 185
rect -210 154 -136 169
rect -546 102 -480 121
rect -546 62 -535 102
rect -495 62 -480 102
rect -210 114 -196 154
rect -151 114 -136 154
rect -26 163 23 168
rect -26 124 -22 163
rect 18 124 23 163
rect 993 153 997 180
rect 1026 153 1031 180
rect 993 149 1031 153
rect 1001 133 1021 149
rect 1150 133 1171 192
rect 3687 188 3694 219
rect 3727 203 3733 219
rect 3727 188 3811 203
rect 3687 182 3811 188
rect 2136 133 3763 163
rect -26 120 23 124
rect 993 125 1031 133
rect -210 99 -136 114
rect 842 96 880 121
rect 993 108 1002 125
rect 1022 108 1031 125
rect 993 101 1031 108
rect 1143 125 1181 133
rect 1143 108 1152 125
rect 1172 108 1181 125
rect 1143 101 1181 108
rect 1978 112 2020 120
rect 2136 112 2162 133
rect 1978 104 2162 112
rect 3729 121 3763 133
rect -546 51 -480 62
rect 42 74 78 79
rect 42 42 47 74
rect 73 42 78 74
rect -227 31 -176 41
rect -227 -2 -221 31
rect -181 -2 -176 31
rect 42 28 51 42
rect 69 28 78 42
rect 842 78 850 96
rect 868 78 880 96
rect 842 61 880 78
rect 1978 86 1991 104
rect 2009 86 2162 104
rect 1978 85 2162 86
rect 2192 100 2250 108
rect 1978 75 2020 85
rect 2192 83 2225 100
rect 2243 83 2250 100
rect 2192 77 2250 83
rect 3729 103 3735 121
rect 3753 103 3763 121
rect 3729 84 3763 103
rect 2192 61 2220 77
rect 42 20 78 28
rect 553 28 622 37
rect 842 34 2220 61
rect 3729 66 3735 84
rect 3753 66 3763 84
rect 3729 39 3763 66
rect 3788 78 3811 182
rect 5223 125 5259 129
rect 5223 99 5226 125
rect 5255 99 5259 125
rect 5223 90 5259 99
rect 3788 70 3836 78
rect 3788 42 3794 70
rect 3830 42 3836 70
rect 5229 49 5253 90
rect 3788 35 3836 42
rect 5224 41 5257 49
rect -227 -7 -176 -2
rect 553 0 565 28
rect 614 0 622 28
rect 5224 23 5232 41
rect 5250 23 5257 41
rect 5224 14 5257 23
rect 553 -6 622 0
<< via1 >>
rect -499 643 -450 646
rect -499 620 -489 643
rect -489 620 -464 643
rect -464 620 -450 643
rect -499 615 -450 620
rect 1218 642 1282 647
rect 1218 620 1236 642
rect 1236 620 1262 642
rect 1262 620 1282 642
rect 1218 609 1282 620
rect 2834 644 2891 645
rect 2834 618 2849 644
rect 2849 618 2876 644
rect 2876 618 2891 644
rect 2834 613 2891 618
rect 1157 431 1197 467
rect -660 317 -618 323
rect -660 296 -651 317
rect -651 296 -627 317
rect -627 296 -618 317
rect -660 289 -618 296
rect -409 319 -372 327
rect -409 296 -403 319
rect -403 296 -379 319
rect -379 296 -372 319
rect -409 288 -372 296
rect 4354 644 4395 649
rect 4354 621 4361 644
rect 4361 621 4387 644
rect 4387 621 4395 644
rect 4354 617 4395 621
rect -535 62 -495 102
rect -196 114 -151 154
rect -22 153 18 163
rect -22 134 -12 153
rect -12 134 7 153
rect 7 134 18 153
rect -22 124 18 134
rect 997 153 1026 180
rect 3694 215 3727 219
rect 3694 192 3699 215
rect 3699 192 3721 215
rect 3721 192 3727 215
rect 3694 188 3727 192
rect 47 46 73 74
rect 47 42 51 46
rect 51 42 69 46
rect 69 42 73 46
rect -221 26 -181 31
rect -221 2 -213 26
rect -213 2 -188 26
rect -188 2 -181 26
rect -221 -2 -181 2
rect 5226 99 5255 125
rect 3794 42 3830 70
rect 565 19 614 28
rect 565 1 578 19
rect 578 1 598 19
rect 598 1 614 19
rect 565 0 614 1
<< metal2 >>
rect -694 649 5271 653
rect -694 647 4354 649
rect -694 646 1218 647
rect -694 625 -499 646
rect -508 615 -499 625
rect -450 625 1218 646
rect -450 615 -444 625
rect -19 623 552 625
rect -508 609 -444 615
rect 1206 609 1218 625
rect 1282 645 4354 647
rect 1282 625 2834 645
rect 1282 609 1294 625
rect 1206 603 1294 609
rect 2826 613 2834 625
rect 2891 625 4354 645
rect 2891 613 2899 625
rect 2826 607 2899 613
rect 4348 617 4354 625
rect 4395 625 5271 649
rect 4395 617 4400 625
rect 4348 611 4400 617
rect 1151 467 1203 473
rect 1151 431 1157 467
rect 1197 462 1203 467
rect 1197 433 5271 462
rect 1197 431 1203 433
rect 1151 425 1203 431
rect 2619 387 5271 411
rect 2619 376 2641 387
rect -702 353 2641 376
rect -670 323 -609 330
rect -670 322 -660 323
rect -701 294 -660 322
rect -670 289 -660 294
rect -618 289 -609 323
rect -670 283 -609 289
rect -419 327 -364 333
rect -419 288 -409 327
rect -372 288 -364 327
rect -419 282 -364 288
rect -401 264 -375 282
rect -699 236 -375 264
rect 3647 242 5250 262
rect 3686 219 3734 226
rect -702 192 1020 215
rect 993 185 1020 192
rect 3686 188 3694 219
rect 3727 188 3734 219
rect 993 180 1031 185
rect 3686 182 3734 188
rect -210 154 -136 169
rect -546 102 -480 121
rect -546 62 -535 102
rect -495 80 -480 102
rect -210 114 -196 154
rect -151 150 -136 154
rect -26 163 34 168
rect -26 151 -22 163
rect -86 150 -22 151
rect -151 124 -22 150
rect 18 124 34 163
rect 993 153 997 180
rect 1026 153 1031 180
rect 993 149 1031 153
rect 5223 125 5259 129
rect -151 122 5122 124
rect 5223 122 5226 125
rect -151 119 5226 122
rect -151 117 -66 119
rect -151 114 -136 117
rect -210 99 -136 114
rect 10 99 5226 119
rect 5255 122 5259 125
rect 5255 99 5271 122
rect 10 98 5271 99
rect 10 95 5122 98
rect 5223 94 5259 98
rect -495 79 -44 80
rect -495 74 5271 79
rect -495 62 47 74
rect -546 51 47 62
rect 42 42 47 51
rect 73 70 5271 74
rect 73 59 3794 70
rect 73 42 78 59
rect -227 31 -176 37
rect 42 36 78 42
rect 3788 42 3794 59
rect 3830 59 5271 70
rect 3830 42 3836 59
rect -227 17 -221 31
rect -671 -2 -221 17
rect -181 17 -176 31
rect 553 28 622 37
rect 3788 35 3836 42
rect 553 17 565 28
rect -181 0 565 17
rect 614 17 622 28
rect 614 0 5267 17
rect -181 -2 5267 0
rect -671 -6 5267 -2
rect -227 -7 -176 -6
<< end >>
