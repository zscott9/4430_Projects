* Diff Pair Bias Trans
X0 nint pbias vdd vdd sky130_fd_pr__pfet_01v8 w=6.0 l=0.4
* Diff In +
X1 n14 vin1 nint vdd sky130_fd_pr__pfet_01v8 w=18 l=1.0
* Diff in -
X2 n23 vin2 nint vdd sky130_fd_pr__pfet_01v8 w=18 l=1.0
* Bias Trans 1
X3 n14 nbias gnd gnd sky130_fd_pr__nfet_01v8 w=6 l=2.0
* Bias Trans 2
X4 n23 nbias gnd gnd sky130_fd_pr__nfet_01v8 w=6 l=2.0
* B1 nFET1
X5 n810 ncasc n14 gnd sky130_fd_pr__nfet_01v8 w=3.0 l=2.0
* B1 pFET1
X6 n810 pcasc n68 vdd sky130_fd_pr__pfet_01v8 w=3.0 l=2.0
* B1 pFET2
X7 n68 n810 vdd vdd sky130_fd_pr__pfet_01v8 w=3.0 l=2.0
* B2 nFET1
X8 n79 ncasc n23 gnd sky130_fd_pr__nfet_01v8 w=3.0 l=2.0
* B2 pFET1
X9 n79 pcasc n57 vdd sky130_fd_pr__pfet_01v8 w=3.0 l=2.0
* B2 pFET2
X10 n57 n810 vdd vdd sky130_fd_pr__pfet_01v8 w=3.0 l=2.0
* Circuit to Set P-Cascode Gate Voltages
X11 psc psc vdd vdd sky130_fd_pr__pfet_01v8 w=3 l=2
X12 pcasc pcasc psc vdd sky130_fd_pr__pfet_01v8 w=3 l=2
X13 pcasc nbias gnd gnd sky130_fd_pr__nfet_01v8 w=0.8 l=0.4
* Circuit to Set N-Cascode Gate Voltages
X14 ncasc ncasc nsc gnd sky130_fd_pr__nfet_01v8 w=3 l=2
X15 nsc nsc gnd gnd sky130_fd_pr__nfet_01v8 w=3 l=2
X16 ncasc pbias vdd vdd sky130_fd_pr__pfet_01v8 w=0.8 l=0.4